module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  wire [63:0] _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  wire [63:0] _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  wire [63:0] _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  wire [63:0] _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  wire [63:0] _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT(
  input         clock,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_8_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_8_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_8_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_9_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_9_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_9_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_10_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_10_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_10_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_10_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_10_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [11:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [11:0] _T_1 = cnt + 12'h1; // @[FFT.scala 42:16]
  reg [11:0] cntD1; // @[FFT.scala 44:22]
  reg [31:0] _RAND_1;
  wire [31:0] _GEN_4 = 11'h3 == cnt[10:0] ? $signed(32'shffff) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_5 = 11'h4 == cnt[10:0] ? $signed(32'shffff) : $signed(_GEN_4); // @[FFT.scala 34:12]
  wire [31:0] _GEN_6 = 11'h5 == cnt[10:0] ? $signed(32'shfffe) : $signed(_GEN_5); // @[FFT.scala 34:12]
  wire [31:0] _GEN_7 = 11'h6 == cnt[10:0] ? $signed(32'shfffd) : $signed(_GEN_6); // @[FFT.scala 34:12]
  wire [31:0] _GEN_8 = 11'h7 == cnt[10:0] ? $signed(32'shfffc) : $signed(_GEN_7); // @[FFT.scala 34:12]
  wire [31:0] _GEN_9 = 11'h8 == cnt[10:0] ? $signed(32'shfffb) : $signed(_GEN_8); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10 = 11'h9 == cnt[10:0] ? $signed(32'shfffa) : $signed(_GEN_9); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11 = 11'ha == cnt[10:0] ? $signed(32'shfff8) : $signed(_GEN_10); // @[FFT.scala 34:12]
  wire [31:0] _GEN_12 = 11'hb == cnt[10:0] ? $signed(32'shfff7) : $signed(_GEN_11); // @[FFT.scala 34:12]
  wire [31:0] _GEN_13 = 11'hc == cnt[10:0] ? $signed(32'shfff5) : $signed(_GEN_12); // @[FFT.scala 34:12]
  wire [31:0] _GEN_14 = 11'hd == cnt[10:0] ? $signed(32'shfff3) : $signed(_GEN_13); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15 = 11'he == cnt[10:0] ? $signed(32'shfff1) : $signed(_GEN_14); // @[FFT.scala 34:12]
  wire [31:0] _GEN_16 = 11'hf == cnt[10:0] ? $signed(32'shffef) : $signed(_GEN_15); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17 = 11'h10 == cnt[10:0] ? $signed(32'shffec) : $signed(_GEN_16); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18 = 11'h11 == cnt[10:0] ? $signed(32'shffea) : $signed(_GEN_17); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19 = 11'h12 == cnt[10:0] ? $signed(32'shffe7) : $signed(_GEN_18); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20 = 11'h13 == cnt[10:0] ? $signed(32'shffe4) : $signed(_GEN_19); // @[FFT.scala 34:12]
  wire [31:0] _GEN_21 = 11'h14 == cnt[10:0] ? $signed(32'shffe1) : $signed(_GEN_20); // @[FFT.scala 34:12]
  wire [31:0] _GEN_22 = 11'h15 == cnt[10:0] ? $signed(32'shffde) : $signed(_GEN_21); // @[FFT.scala 34:12]
  wire [31:0] _GEN_23 = 11'h16 == cnt[10:0] ? $signed(32'shffdb) : $signed(_GEN_22); // @[FFT.scala 34:12]
  wire [31:0] _GEN_24 = 11'h17 == cnt[10:0] ? $signed(32'shffd7) : $signed(_GEN_23); // @[FFT.scala 34:12]
  wire [31:0] _GEN_25 = 11'h18 == cnt[10:0] ? $signed(32'shffd4) : $signed(_GEN_24); // @[FFT.scala 34:12]
  wire [31:0] _GEN_26 = 11'h19 == cnt[10:0] ? $signed(32'shffd0) : $signed(_GEN_25); // @[FFT.scala 34:12]
  wire [31:0] _GEN_27 = 11'h1a == cnt[10:0] ? $signed(32'shffcc) : $signed(_GEN_26); // @[FFT.scala 34:12]
  wire [31:0] _GEN_28 = 11'h1b == cnt[10:0] ? $signed(32'shffc8) : $signed(_GEN_27); // @[FFT.scala 34:12]
  wire [31:0] _GEN_29 = 11'h1c == cnt[10:0] ? $signed(32'shffc4) : $signed(_GEN_28); // @[FFT.scala 34:12]
  wire [31:0] _GEN_30 = 11'h1d == cnt[10:0] ? $signed(32'shffbf) : $signed(_GEN_29); // @[FFT.scala 34:12]
  wire [31:0] _GEN_31 = 11'h1e == cnt[10:0] ? $signed(32'shffbb) : $signed(_GEN_30); // @[FFT.scala 34:12]
  wire [31:0] _GEN_32 = 11'h1f == cnt[10:0] ? $signed(32'shffb6) : $signed(_GEN_31); // @[FFT.scala 34:12]
  wire [31:0] _GEN_33 = 11'h20 == cnt[10:0] ? $signed(32'shffb1) : $signed(_GEN_32); // @[FFT.scala 34:12]
  wire [31:0] _GEN_34 = 11'h21 == cnt[10:0] ? $signed(32'shffac) : $signed(_GEN_33); // @[FFT.scala 34:12]
  wire [31:0] _GEN_35 = 11'h22 == cnt[10:0] ? $signed(32'shffa7) : $signed(_GEN_34); // @[FFT.scala 34:12]
  wire [31:0] _GEN_36 = 11'h23 == cnt[10:0] ? $signed(32'shffa2) : $signed(_GEN_35); // @[FFT.scala 34:12]
  wire [31:0] _GEN_37 = 11'h24 == cnt[10:0] ? $signed(32'shff9c) : $signed(_GEN_36); // @[FFT.scala 34:12]
  wire [31:0] _GEN_38 = 11'h25 == cnt[10:0] ? $signed(32'shff96) : $signed(_GEN_37); // @[FFT.scala 34:12]
  wire [31:0] _GEN_39 = 11'h26 == cnt[10:0] ? $signed(32'shff91) : $signed(_GEN_38); // @[FFT.scala 34:12]
  wire [31:0] _GEN_40 = 11'h27 == cnt[10:0] ? $signed(32'shff8b) : $signed(_GEN_39); // @[FFT.scala 34:12]
  wire [31:0] _GEN_41 = 11'h28 == cnt[10:0] ? $signed(32'shff85) : $signed(_GEN_40); // @[FFT.scala 34:12]
  wire [31:0] _GEN_42 = 11'h29 == cnt[10:0] ? $signed(32'shff7e) : $signed(_GEN_41); // @[FFT.scala 34:12]
  wire [31:0] _GEN_43 = 11'h2a == cnt[10:0] ? $signed(32'shff78) : $signed(_GEN_42); // @[FFT.scala 34:12]
  wire [31:0] _GEN_44 = 11'h2b == cnt[10:0] ? $signed(32'shff71) : $signed(_GEN_43); // @[FFT.scala 34:12]
  wire [31:0] _GEN_45 = 11'h2c == cnt[10:0] ? $signed(32'shff6b) : $signed(_GEN_44); // @[FFT.scala 34:12]
  wire [31:0] _GEN_46 = 11'h2d == cnt[10:0] ? $signed(32'shff64) : $signed(_GEN_45); // @[FFT.scala 34:12]
  wire [31:0] _GEN_47 = 11'h2e == cnt[10:0] ? $signed(32'shff5d) : $signed(_GEN_46); // @[FFT.scala 34:12]
  wire [31:0] _GEN_48 = 11'h2f == cnt[10:0] ? $signed(32'shff56) : $signed(_GEN_47); // @[FFT.scala 34:12]
  wire [31:0] _GEN_49 = 11'h30 == cnt[10:0] ? $signed(32'shff4e) : $signed(_GEN_48); // @[FFT.scala 34:12]
  wire [31:0] _GEN_50 = 11'h31 == cnt[10:0] ? $signed(32'shff47) : $signed(_GEN_49); // @[FFT.scala 34:12]
  wire [31:0] _GEN_51 = 11'h32 == cnt[10:0] ? $signed(32'shff3f) : $signed(_GEN_50); // @[FFT.scala 34:12]
  wire [31:0] _GEN_52 = 11'h33 == cnt[10:0] ? $signed(32'shff38) : $signed(_GEN_51); // @[FFT.scala 34:12]
  wire [31:0] _GEN_53 = 11'h34 == cnt[10:0] ? $signed(32'shff30) : $signed(_GEN_52); // @[FFT.scala 34:12]
  wire [31:0] _GEN_54 = 11'h35 == cnt[10:0] ? $signed(32'shff28) : $signed(_GEN_53); // @[FFT.scala 34:12]
  wire [31:0] _GEN_55 = 11'h36 == cnt[10:0] ? $signed(32'shff1f) : $signed(_GEN_54); // @[FFT.scala 34:12]
  wire [31:0] _GEN_56 = 11'h37 == cnt[10:0] ? $signed(32'shff17) : $signed(_GEN_55); // @[FFT.scala 34:12]
  wire [31:0] _GEN_57 = 11'h38 == cnt[10:0] ? $signed(32'shff0e) : $signed(_GEN_56); // @[FFT.scala 34:12]
  wire [31:0] _GEN_58 = 11'h39 == cnt[10:0] ? $signed(32'shff06) : $signed(_GEN_57); // @[FFT.scala 34:12]
  wire [31:0] _GEN_59 = 11'h3a == cnt[10:0] ? $signed(32'shfefd) : $signed(_GEN_58); // @[FFT.scala 34:12]
  wire [31:0] _GEN_60 = 11'h3b == cnt[10:0] ? $signed(32'shfef4) : $signed(_GEN_59); // @[FFT.scala 34:12]
  wire [31:0] _GEN_61 = 11'h3c == cnt[10:0] ? $signed(32'shfeeb) : $signed(_GEN_60); // @[FFT.scala 34:12]
  wire [31:0] _GEN_62 = 11'h3d == cnt[10:0] ? $signed(32'shfee1) : $signed(_GEN_61); // @[FFT.scala 34:12]
  wire [31:0] _GEN_63 = 11'h3e == cnt[10:0] ? $signed(32'shfed8) : $signed(_GEN_62); // @[FFT.scala 34:12]
  wire [31:0] _GEN_64 = 11'h3f == cnt[10:0] ? $signed(32'shfece) : $signed(_GEN_63); // @[FFT.scala 34:12]
  wire [31:0] _GEN_65 = 11'h40 == cnt[10:0] ? $signed(32'shfec4) : $signed(_GEN_64); // @[FFT.scala 34:12]
  wire [31:0] _GEN_66 = 11'h41 == cnt[10:0] ? $signed(32'shfeba) : $signed(_GEN_65); // @[FFT.scala 34:12]
  wire [31:0] _GEN_67 = 11'h42 == cnt[10:0] ? $signed(32'shfeb0) : $signed(_GEN_66); // @[FFT.scala 34:12]
  wire [31:0] _GEN_68 = 11'h43 == cnt[10:0] ? $signed(32'shfea6) : $signed(_GEN_67); // @[FFT.scala 34:12]
  wire [31:0] _GEN_69 = 11'h44 == cnt[10:0] ? $signed(32'shfe9c) : $signed(_GEN_68); // @[FFT.scala 34:12]
  wire [31:0] _GEN_70 = 11'h45 == cnt[10:0] ? $signed(32'shfe91) : $signed(_GEN_69); // @[FFT.scala 34:12]
  wire [31:0] _GEN_71 = 11'h46 == cnt[10:0] ? $signed(32'shfe87) : $signed(_GEN_70); // @[FFT.scala 34:12]
  wire [31:0] _GEN_72 = 11'h47 == cnt[10:0] ? $signed(32'shfe7c) : $signed(_GEN_71); // @[FFT.scala 34:12]
  wire [31:0] _GEN_73 = 11'h48 == cnt[10:0] ? $signed(32'shfe71) : $signed(_GEN_72); // @[FFT.scala 34:12]
  wire [31:0] _GEN_74 = 11'h49 == cnt[10:0] ? $signed(32'shfe66) : $signed(_GEN_73); // @[FFT.scala 34:12]
  wire [31:0] _GEN_75 = 11'h4a == cnt[10:0] ? $signed(32'shfe5a) : $signed(_GEN_74); // @[FFT.scala 34:12]
  wire [31:0] _GEN_76 = 11'h4b == cnt[10:0] ? $signed(32'shfe4f) : $signed(_GEN_75); // @[FFT.scala 34:12]
  wire [31:0] _GEN_77 = 11'h4c == cnt[10:0] ? $signed(32'shfe43) : $signed(_GEN_76); // @[FFT.scala 34:12]
  wire [31:0] _GEN_78 = 11'h4d == cnt[10:0] ? $signed(32'shfe37) : $signed(_GEN_77); // @[FFT.scala 34:12]
  wire [31:0] _GEN_79 = 11'h4e == cnt[10:0] ? $signed(32'shfe2b) : $signed(_GEN_78); // @[FFT.scala 34:12]
  wire [31:0] _GEN_80 = 11'h4f == cnt[10:0] ? $signed(32'shfe1f) : $signed(_GEN_79); // @[FFT.scala 34:12]
  wire [31:0] _GEN_81 = 11'h50 == cnt[10:0] ? $signed(32'shfe13) : $signed(_GEN_80); // @[FFT.scala 34:12]
  wire [31:0] _GEN_82 = 11'h51 == cnt[10:0] ? $signed(32'shfe07) : $signed(_GEN_81); // @[FFT.scala 34:12]
  wire [31:0] _GEN_83 = 11'h52 == cnt[10:0] ? $signed(32'shfdfa) : $signed(_GEN_82); // @[FFT.scala 34:12]
  wire [31:0] _GEN_84 = 11'h53 == cnt[10:0] ? $signed(32'shfdee) : $signed(_GEN_83); // @[FFT.scala 34:12]
  wire [31:0] _GEN_85 = 11'h54 == cnt[10:0] ? $signed(32'shfde1) : $signed(_GEN_84); // @[FFT.scala 34:12]
  wire [31:0] _GEN_86 = 11'h55 == cnt[10:0] ? $signed(32'shfdd4) : $signed(_GEN_85); // @[FFT.scala 34:12]
  wire [31:0] _GEN_87 = 11'h56 == cnt[10:0] ? $signed(32'shfdc7) : $signed(_GEN_86); // @[FFT.scala 34:12]
  wire [31:0] _GEN_88 = 11'h57 == cnt[10:0] ? $signed(32'shfdb9) : $signed(_GEN_87); // @[FFT.scala 34:12]
  wire [31:0] _GEN_89 = 11'h58 == cnt[10:0] ? $signed(32'shfdac) : $signed(_GEN_88); // @[FFT.scala 34:12]
  wire [31:0] _GEN_90 = 11'h59 == cnt[10:0] ? $signed(32'shfd9e) : $signed(_GEN_89); // @[FFT.scala 34:12]
  wire [31:0] _GEN_91 = 11'h5a == cnt[10:0] ? $signed(32'shfd90) : $signed(_GEN_90); // @[FFT.scala 34:12]
  wire [31:0] _GEN_92 = 11'h5b == cnt[10:0] ? $signed(32'shfd83) : $signed(_GEN_91); // @[FFT.scala 34:12]
  wire [31:0] _GEN_93 = 11'h5c == cnt[10:0] ? $signed(32'shfd74) : $signed(_GEN_92); // @[FFT.scala 34:12]
  wire [31:0] _GEN_94 = 11'h5d == cnt[10:0] ? $signed(32'shfd66) : $signed(_GEN_93); // @[FFT.scala 34:12]
  wire [31:0] _GEN_95 = 11'h5e == cnt[10:0] ? $signed(32'shfd58) : $signed(_GEN_94); // @[FFT.scala 34:12]
  wire [31:0] _GEN_96 = 11'h5f == cnt[10:0] ? $signed(32'shfd49) : $signed(_GEN_95); // @[FFT.scala 34:12]
  wire [31:0] _GEN_97 = 11'h60 == cnt[10:0] ? $signed(32'shfd3b) : $signed(_GEN_96); // @[FFT.scala 34:12]
  wire [31:0] _GEN_98 = 11'h61 == cnt[10:0] ? $signed(32'shfd2c) : $signed(_GEN_97); // @[FFT.scala 34:12]
  wire [31:0] _GEN_99 = 11'h62 == cnt[10:0] ? $signed(32'shfd1d) : $signed(_GEN_98); // @[FFT.scala 34:12]
  wire [31:0] _GEN_100 = 11'h63 == cnt[10:0] ? $signed(32'shfd0e) : $signed(_GEN_99); // @[FFT.scala 34:12]
  wire [31:0] _GEN_101 = 11'h64 == cnt[10:0] ? $signed(32'shfcfe) : $signed(_GEN_100); // @[FFT.scala 34:12]
  wire [31:0] _GEN_102 = 11'h65 == cnt[10:0] ? $signed(32'shfcef) : $signed(_GEN_101); // @[FFT.scala 34:12]
  wire [31:0] _GEN_103 = 11'h66 == cnt[10:0] ? $signed(32'shfcdf) : $signed(_GEN_102); // @[FFT.scala 34:12]
  wire [31:0] _GEN_104 = 11'h67 == cnt[10:0] ? $signed(32'shfcd0) : $signed(_GEN_103); // @[FFT.scala 34:12]
  wire [31:0] _GEN_105 = 11'h68 == cnt[10:0] ? $signed(32'shfcc0) : $signed(_GEN_104); // @[FFT.scala 34:12]
  wire [31:0] _GEN_106 = 11'h69 == cnt[10:0] ? $signed(32'shfcb0) : $signed(_GEN_105); // @[FFT.scala 34:12]
  wire [31:0] _GEN_107 = 11'h6a == cnt[10:0] ? $signed(32'shfca0) : $signed(_GEN_106); // @[FFT.scala 34:12]
  wire [31:0] _GEN_108 = 11'h6b == cnt[10:0] ? $signed(32'shfc8f) : $signed(_GEN_107); // @[FFT.scala 34:12]
  wire [31:0] _GEN_109 = 11'h6c == cnt[10:0] ? $signed(32'shfc7f) : $signed(_GEN_108); // @[FFT.scala 34:12]
  wire [31:0] _GEN_110 = 11'h6d == cnt[10:0] ? $signed(32'shfc6e) : $signed(_GEN_109); // @[FFT.scala 34:12]
  wire [31:0] _GEN_111 = 11'h6e == cnt[10:0] ? $signed(32'shfc5d) : $signed(_GEN_110); // @[FFT.scala 34:12]
  wire [31:0] _GEN_112 = 11'h6f == cnt[10:0] ? $signed(32'shfc4c) : $signed(_GEN_111); // @[FFT.scala 34:12]
  wire [31:0] _GEN_113 = 11'h70 == cnt[10:0] ? $signed(32'shfc3b) : $signed(_GEN_112); // @[FFT.scala 34:12]
  wire [31:0] _GEN_114 = 11'h71 == cnt[10:0] ? $signed(32'shfc2a) : $signed(_GEN_113); // @[FFT.scala 34:12]
  wire [31:0] _GEN_115 = 11'h72 == cnt[10:0] ? $signed(32'shfc18) : $signed(_GEN_114); // @[FFT.scala 34:12]
  wire [31:0] _GEN_116 = 11'h73 == cnt[10:0] ? $signed(32'shfc07) : $signed(_GEN_115); // @[FFT.scala 34:12]
  wire [31:0] _GEN_117 = 11'h74 == cnt[10:0] ? $signed(32'shfbf5) : $signed(_GEN_116); // @[FFT.scala 34:12]
  wire [31:0] _GEN_118 = 11'h75 == cnt[10:0] ? $signed(32'shfbe3) : $signed(_GEN_117); // @[FFT.scala 34:12]
  wire [31:0] _GEN_119 = 11'h76 == cnt[10:0] ? $signed(32'shfbd1) : $signed(_GEN_118); // @[FFT.scala 34:12]
  wire [31:0] _GEN_120 = 11'h77 == cnt[10:0] ? $signed(32'shfbbf) : $signed(_GEN_119); // @[FFT.scala 34:12]
  wire [31:0] _GEN_121 = 11'h78 == cnt[10:0] ? $signed(32'shfbad) : $signed(_GEN_120); // @[FFT.scala 34:12]
  wire [31:0] _GEN_122 = 11'h79 == cnt[10:0] ? $signed(32'shfb9a) : $signed(_GEN_121); // @[FFT.scala 34:12]
  wire [31:0] _GEN_123 = 11'h7a == cnt[10:0] ? $signed(32'shfb88) : $signed(_GEN_122); // @[FFT.scala 34:12]
  wire [31:0] _GEN_124 = 11'h7b == cnt[10:0] ? $signed(32'shfb75) : $signed(_GEN_123); // @[FFT.scala 34:12]
  wire [31:0] _GEN_125 = 11'h7c == cnt[10:0] ? $signed(32'shfb62) : $signed(_GEN_124); // @[FFT.scala 34:12]
  wire [31:0] _GEN_126 = 11'h7d == cnt[10:0] ? $signed(32'shfb4f) : $signed(_GEN_125); // @[FFT.scala 34:12]
  wire [31:0] _GEN_127 = 11'h7e == cnt[10:0] ? $signed(32'shfb3c) : $signed(_GEN_126); // @[FFT.scala 34:12]
  wire [31:0] _GEN_128 = 11'h7f == cnt[10:0] ? $signed(32'shfb28) : $signed(_GEN_127); // @[FFT.scala 34:12]
  wire [31:0] _GEN_129 = 11'h80 == cnt[10:0] ? $signed(32'shfb15) : $signed(_GEN_128); // @[FFT.scala 34:12]
  wire [31:0] _GEN_130 = 11'h81 == cnt[10:0] ? $signed(32'shfb01) : $signed(_GEN_129); // @[FFT.scala 34:12]
  wire [31:0] _GEN_131 = 11'h82 == cnt[10:0] ? $signed(32'shfaed) : $signed(_GEN_130); // @[FFT.scala 34:12]
  wire [31:0] _GEN_132 = 11'h83 == cnt[10:0] ? $signed(32'shfad9) : $signed(_GEN_131); // @[FFT.scala 34:12]
  wire [31:0] _GEN_133 = 11'h84 == cnt[10:0] ? $signed(32'shfac5) : $signed(_GEN_132); // @[FFT.scala 34:12]
  wire [31:0] _GEN_134 = 11'h85 == cnt[10:0] ? $signed(32'shfab1) : $signed(_GEN_133); // @[FFT.scala 34:12]
  wire [31:0] _GEN_135 = 11'h86 == cnt[10:0] ? $signed(32'shfa9c) : $signed(_GEN_134); // @[FFT.scala 34:12]
  wire [31:0] _GEN_136 = 11'h87 == cnt[10:0] ? $signed(32'shfa88) : $signed(_GEN_135); // @[FFT.scala 34:12]
  wire [31:0] _GEN_137 = 11'h88 == cnt[10:0] ? $signed(32'shfa73) : $signed(_GEN_136); // @[FFT.scala 34:12]
  wire [31:0] _GEN_138 = 11'h89 == cnt[10:0] ? $signed(32'shfa5e) : $signed(_GEN_137); // @[FFT.scala 34:12]
  wire [31:0] _GEN_139 = 11'h8a == cnt[10:0] ? $signed(32'shfa49) : $signed(_GEN_138); // @[FFT.scala 34:12]
  wire [31:0] _GEN_140 = 11'h8b == cnt[10:0] ? $signed(32'shfa34) : $signed(_GEN_139); // @[FFT.scala 34:12]
  wire [31:0] _GEN_141 = 11'h8c == cnt[10:0] ? $signed(32'shfa1f) : $signed(_GEN_140); // @[FFT.scala 34:12]
  wire [31:0] _GEN_142 = 11'h8d == cnt[10:0] ? $signed(32'shfa09) : $signed(_GEN_141); // @[FFT.scala 34:12]
  wire [31:0] _GEN_143 = 11'h8e == cnt[10:0] ? $signed(32'shf9f3) : $signed(_GEN_142); // @[FFT.scala 34:12]
  wire [31:0] _GEN_144 = 11'h8f == cnt[10:0] ? $signed(32'shf9de) : $signed(_GEN_143); // @[FFT.scala 34:12]
  wire [31:0] _GEN_145 = 11'h90 == cnt[10:0] ? $signed(32'shf9c8) : $signed(_GEN_144); // @[FFT.scala 34:12]
  wire [31:0] _GEN_146 = 11'h91 == cnt[10:0] ? $signed(32'shf9b2) : $signed(_GEN_145); // @[FFT.scala 34:12]
  wire [31:0] _GEN_147 = 11'h92 == cnt[10:0] ? $signed(32'shf99b) : $signed(_GEN_146); // @[FFT.scala 34:12]
  wire [31:0] _GEN_148 = 11'h93 == cnt[10:0] ? $signed(32'shf985) : $signed(_GEN_147); // @[FFT.scala 34:12]
  wire [31:0] _GEN_149 = 11'h94 == cnt[10:0] ? $signed(32'shf96e) : $signed(_GEN_148); // @[FFT.scala 34:12]
  wire [31:0] _GEN_150 = 11'h95 == cnt[10:0] ? $signed(32'shf958) : $signed(_GEN_149); // @[FFT.scala 34:12]
  wire [31:0] _GEN_151 = 11'h96 == cnt[10:0] ? $signed(32'shf941) : $signed(_GEN_150); // @[FFT.scala 34:12]
  wire [31:0] _GEN_152 = 11'h97 == cnt[10:0] ? $signed(32'shf92a) : $signed(_GEN_151); // @[FFT.scala 34:12]
  wire [31:0] _GEN_153 = 11'h98 == cnt[10:0] ? $signed(32'shf913) : $signed(_GEN_152); // @[FFT.scala 34:12]
  wire [31:0] _GEN_154 = 11'h99 == cnt[10:0] ? $signed(32'shf8fb) : $signed(_GEN_153); // @[FFT.scala 34:12]
  wire [31:0] _GEN_155 = 11'h9a == cnt[10:0] ? $signed(32'shf8e4) : $signed(_GEN_154); // @[FFT.scala 34:12]
  wire [31:0] _GEN_156 = 11'h9b == cnt[10:0] ? $signed(32'shf8cc) : $signed(_GEN_155); // @[FFT.scala 34:12]
  wire [31:0] _GEN_157 = 11'h9c == cnt[10:0] ? $signed(32'shf8b4) : $signed(_GEN_156); // @[FFT.scala 34:12]
  wire [31:0] _GEN_158 = 11'h9d == cnt[10:0] ? $signed(32'shf89d) : $signed(_GEN_157); // @[FFT.scala 34:12]
  wire [31:0] _GEN_159 = 11'h9e == cnt[10:0] ? $signed(32'shf885) : $signed(_GEN_158); // @[FFT.scala 34:12]
  wire [31:0] _GEN_160 = 11'h9f == cnt[10:0] ? $signed(32'shf86c) : $signed(_GEN_159); // @[FFT.scala 34:12]
  wire [31:0] _GEN_161 = 11'ha0 == cnt[10:0] ? $signed(32'shf854) : $signed(_GEN_160); // @[FFT.scala 34:12]
  wire [31:0] _GEN_162 = 11'ha1 == cnt[10:0] ? $signed(32'shf83b) : $signed(_GEN_161); // @[FFT.scala 34:12]
  wire [31:0] _GEN_163 = 11'ha2 == cnt[10:0] ? $signed(32'shf823) : $signed(_GEN_162); // @[FFT.scala 34:12]
  wire [31:0] _GEN_164 = 11'ha3 == cnt[10:0] ? $signed(32'shf80a) : $signed(_GEN_163); // @[FFT.scala 34:12]
  wire [31:0] _GEN_165 = 11'ha4 == cnt[10:0] ? $signed(32'shf7f1) : $signed(_GEN_164); // @[FFT.scala 34:12]
  wire [31:0] _GEN_166 = 11'ha5 == cnt[10:0] ? $signed(32'shf7d8) : $signed(_GEN_165); // @[FFT.scala 34:12]
  wire [31:0] _GEN_167 = 11'ha6 == cnt[10:0] ? $signed(32'shf7bf) : $signed(_GEN_166); // @[FFT.scala 34:12]
  wire [31:0] _GEN_168 = 11'ha7 == cnt[10:0] ? $signed(32'shf7a5) : $signed(_GEN_167); // @[FFT.scala 34:12]
  wire [31:0] _GEN_169 = 11'ha8 == cnt[10:0] ? $signed(32'shf78c) : $signed(_GEN_168); // @[FFT.scala 34:12]
  wire [31:0] _GEN_170 = 11'ha9 == cnt[10:0] ? $signed(32'shf772) : $signed(_GEN_169); // @[FFT.scala 34:12]
  wire [31:0] _GEN_171 = 11'haa == cnt[10:0] ? $signed(32'shf758) : $signed(_GEN_170); // @[FFT.scala 34:12]
  wire [31:0] _GEN_172 = 11'hab == cnt[10:0] ? $signed(32'shf73e) : $signed(_GEN_171); // @[FFT.scala 34:12]
  wire [31:0] _GEN_173 = 11'hac == cnt[10:0] ? $signed(32'shf724) : $signed(_GEN_172); // @[FFT.scala 34:12]
  wire [31:0] _GEN_174 = 11'had == cnt[10:0] ? $signed(32'shf70a) : $signed(_GEN_173); // @[FFT.scala 34:12]
  wire [31:0] _GEN_175 = 11'hae == cnt[10:0] ? $signed(32'shf6ef) : $signed(_GEN_174); // @[FFT.scala 34:12]
  wire [31:0] _GEN_176 = 11'haf == cnt[10:0] ? $signed(32'shf6d5) : $signed(_GEN_175); // @[FFT.scala 34:12]
  wire [31:0] _GEN_177 = 11'hb0 == cnt[10:0] ? $signed(32'shf6ba) : $signed(_GEN_176); // @[FFT.scala 34:12]
  wire [31:0] _GEN_178 = 11'hb1 == cnt[10:0] ? $signed(32'shf69f) : $signed(_GEN_177); // @[FFT.scala 34:12]
  wire [31:0] _GEN_179 = 11'hb2 == cnt[10:0] ? $signed(32'shf684) : $signed(_GEN_178); // @[FFT.scala 34:12]
  wire [31:0] _GEN_180 = 11'hb3 == cnt[10:0] ? $signed(32'shf669) : $signed(_GEN_179); // @[FFT.scala 34:12]
  wire [31:0] _GEN_181 = 11'hb4 == cnt[10:0] ? $signed(32'shf64e) : $signed(_GEN_180); // @[FFT.scala 34:12]
  wire [31:0] _GEN_182 = 11'hb5 == cnt[10:0] ? $signed(32'shf632) : $signed(_GEN_181); // @[FFT.scala 34:12]
  wire [31:0] _GEN_183 = 11'hb6 == cnt[10:0] ? $signed(32'shf616) : $signed(_GEN_182); // @[FFT.scala 34:12]
  wire [31:0] _GEN_184 = 11'hb7 == cnt[10:0] ? $signed(32'shf5fb) : $signed(_GEN_183); // @[FFT.scala 34:12]
  wire [31:0] _GEN_185 = 11'hb8 == cnt[10:0] ? $signed(32'shf5df) : $signed(_GEN_184); // @[FFT.scala 34:12]
  wire [31:0] _GEN_186 = 11'hb9 == cnt[10:0] ? $signed(32'shf5c3) : $signed(_GEN_185); // @[FFT.scala 34:12]
  wire [31:0] _GEN_187 = 11'hba == cnt[10:0] ? $signed(32'shf5a6) : $signed(_GEN_186); // @[FFT.scala 34:12]
  wire [31:0] _GEN_188 = 11'hbb == cnt[10:0] ? $signed(32'shf58a) : $signed(_GEN_187); // @[FFT.scala 34:12]
  wire [31:0] _GEN_189 = 11'hbc == cnt[10:0] ? $signed(32'shf56e) : $signed(_GEN_188); // @[FFT.scala 34:12]
  wire [31:0] _GEN_190 = 11'hbd == cnt[10:0] ? $signed(32'shf551) : $signed(_GEN_189); // @[FFT.scala 34:12]
  wire [31:0] _GEN_191 = 11'hbe == cnt[10:0] ? $signed(32'shf534) : $signed(_GEN_190); // @[FFT.scala 34:12]
  wire [31:0] _GEN_192 = 11'hbf == cnt[10:0] ? $signed(32'shf517) : $signed(_GEN_191); // @[FFT.scala 34:12]
  wire [31:0] _GEN_193 = 11'hc0 == cnt[10:0] ? $signed(32'shf4fa) : $signed(_GEN_192); // @[FFT.scala 34:12]
  wire [31:0] _GEN_194 = 11'hc1 == cnt[10:0] ? $signed(32'shf4dd) : $signed(_GEN_193); // @[FFT.scala 34:12]
  wire [31:0] _GEN_195 = 11'hc2 == cnt[10:0] ? $signed(32'shf4bf) : $signed(_GEN_194); // @[FFT.scala 34:12]
  wire [31:0] _GEN_196 = 11'hc3 == cnt[10:0] ? $signed(32'shf4a2) : $signed(_GEN_195); // @[FFT.scala 34:12]
  wire [31:0] _GEN_197 = 11'hc4 == cnt[10:0] ? $signed(32'shf484) : $signed(_GEN_196); // @[FFT.scala 34:12]
  wire [31:0] _GEN_198 = 11'hc5 == cnt[10:0] ? $signed(32'shf466) : $signed(_GEN_197); // @[FFT.scala 34:12]
  wire [31:0] _GEN_199 = 11'hc6 == cnt[10:0] ? $signed(32'shf448) : $signed(_GEN_198); // @[FFT.scala 34:12]
  wire [31:0] _GEN_200 = 11'hc7 == cnt[10:0] ? $signed(32'shf42a) : $signed(_GEN_199); // @[FFT.scala 34:12]
  wire [31:0] _GEN_201 = 11'hc8 == cnt[10:0] ? $signed(32'shf40c) : $signed(_GEN_200); // @[FFT.scala 34:12]
  wire [31:0] _GEN_202 = 11'hc9 == cnt[10:0] ? $signed(32'shf3ed) : $signed(_GEN_201); // @[FFT.scala 34:12]
  wire [31:0] _GEN_203 = 11'hca == cnt[10:0] ? $signed(32'shf3cf) : $signed(_GEN_202); // @[FFT.scala 34:12]
  wire [31:0] _GEN_204 = 11'hcb == cnt[10:0] ? $signed(32'shf3b0) : $signed(_GEN_203); // @[FFT.scala 34:12]
  wire [31:0] _GEN_205 = 11'hcc == cnt[10:0] ? $signed(32'shf391) : $signed(_GEN_204); // @[FFT.scala 34:12]
  wire [31:0] _GEN_206 = 11'hcd == cnt[10:0] ? $signed(32'shf372) : $signed(_GEN_205); // @[FFT.scala 34:12]
  wire [31:0] _GEN_207 = 11'hce == cnt[10:0] ? $signed(32'shf353) : $signed(_GEN_206); // @[FFT.scala 34:12]
  wire [31:0] _GEN_208 = 11'hcf == cnt[10:0] ? $signed(32'shf334) : $signed(_GEN_207); // @[FFT.scala 34:12]
  wire [31:0] _GEN_209 = 11'hd0 == cnt[10:0] ? $signed(32'shf314) : $signed(_GEN_208); // @[FFT.scala 34:12]
  wire [31:0] _GEN_210 = 11'hd1 == cnt[10:0] ? $signed(32'shf2f5) : $signed(_GEN_209); // @[FFT.scala 34:12]
  wire [31:0] _GEN_211 = 11'hd2 == cnt[10:0] ? $signed(32'shf2d5) : $signed(_GEN_210); // @[FFT.scala 34:12]
  wire [31:0] _GEN_212 = 11'hd3 == cnt[10:0] ? $signed(32'shf2b5) : $signed(_GEN_211); // @[FFT.scala 34:12]
  wire [31:0] _GEN_213 = 11'hd4 == cnt[10:0] ? $signed(32'shf295) : $signed(_GEN_212); // @[FFT.scala 34:12]
  wire [31:0] _GEN_214 = 11'hd5 == cnt[10:0] ? $signed(32'shf275) : $signed(_GEN_213); // @[FFT.scala 34:12]
  wire [31:0] _GEN_215 = 11'hd6 == cnt[10:0] ? $signed(32'shf254) : $signed(_GEN_214); // @[FFT.scala 34:12]
  wire [31:0] _GEN_216 = 11'hd7 == cnt[10:0] ? $signed(32'shf234) : $signed(_GEN_215); // @[FFT.scala 34:12]
  wire [31:0] _GEN_217 = 11'hd8 == cnt[10:0] ? $signed(32'shf213) : $signed(_GEN_216); // @[FFT.scala 34:12]
  wire [31:0] _GEN_218 = 11'hd9 == cnt[10:0] ? $signed(32'shf1f3) : $signed(_GEN_217); // @[FFT.scala 34:12]
  wire [31:0] _GEN_219 = 11'hda == cnt[10:0] ? $signed(32'shf1d2) : $signed(_GEN_218); // @[FFT.scala 34:12]
  wire [31:0] _GEN_220 = 11'hdb == cnt[10:0] ? $signed(32'shf1b1) : $signed(_GEN_219); // @[FFT.scala 34:12]
  wire [31:0] _GEN_221 = 11'hdc == cnt[10:0] ? $signed(32'shf18f) : $signed(_GEN_220); // @[FFT.scala 34:12]
  wire [31:0] _GEN_222 = 11'hdd == cnt[10:0] ? $signed(32'shf16e) : $signed(_GEN_221); // @[FFT.scala 34:12]
  wire [31:0] _GEN_223 = 11'hde == cnt[10:0] ? $signed(32'shf14c) : $signed(_GEN_222); // @[FFT.scala 34:12]
  wire [31:0] _GEN_224 = 11'hdf == cnt[10:0] ? $signed(32'shf12b) : $signed(_GEN_223); // @[FFT.scala 34:12]
  wire [31:0] _GEN_225 = 11'he0 == cnt[10:0] ? $signed(32'shf109) : $signed(_GEN_224); // @[FFT.scala 34:12]
  wire [31:0] _GEN_226 = 11'he1 == cnt[10:0] ? $signed(32'shf0e7) : $signed(_GEN_225); // @[FFT.scala 34:12]
  wire [31:0] _GEN_227 = 11'he2 == cnt[10:0] ? $signed(32'shf0c5) : $signed(_GEN_226); // @[FFT.scala 34:12]
  wire [31:0] _GEN_228 = 11'he3 == cnt[10:0] ? $signed(32'shf0a3) : $signed(_GEN_227); // @[FFT.scala 34:12]
  wire [31:0] _GEN_229 = 11'he4 == cnt[10:0] ? $signed(32'shf080) : $signed(_GEN_228); // @[FFT.scala 34:12]
  wire [31:0] _GEN_230 = 11'he5 == cnt[10:0] ? $signed(32'shf05e) : $signed(_GEN_229); // @[FFT.scala 34:12]
  wire [31:0] _GEN_231 = 11'he6 == cnt[10:0] ? $signed(32'shf03b) : $signed(_GEN_230); // @[FFT.scala 34:12]
  wire [31:0] _GEN_232 = 11'he7 == cnt[10:0] ? $signed(32'shf018) : $signed(_GEN_231); // @[FFT.scala 34:12]
  wire [31:0] _GEN_233 = 11'he8 == cnt[10:0] ? $signed(32'sheff5) : $signed(_GEN_232); // @[FFT.scala 34:12]
  wire [31:0] _GEN_234 = 11'he9 == cnt[10:0] ? $signed(32'shefd2) : $signed(_GEN_233); // @[FFT.scala 34:12]
  wire [31:0] _GEN_235 = 11'hea == cnt[10:0] ? $signed(32'shefaf) : $signed(_GEN_234); // @[FFT.scala 34:12]
  wire [31:0] _GEN_236 = 11'heb == cnt[10:0] ? $signed(32'shef8c) : $signed(_GEN_235); // @[FFT.scala 34:12]
  wire [31:0] _GEN_237 = 11'hec == cnt[10:0] ? $signed(32'shef68) : $signed(_GEN_236); // @[FFT.scala 34:12]
  wire [31:0] _GEN_238 = 11'hed == cnt[10:0] ? $signed(32'shef45) : $signed(_GEN_237); // @[FFT.scala 34:12]
  wire [31:0] _GEN_239 = 11'hee == cnt[10:0] ? $signed(32'shef21) : $signed(_GEN_238); // @[FFT.scala 34:12]
  wire [31:0] _GEN_240 = 11'hef == cnt[10:0] ? $signed(32'sheefd) : $signed(_GEN_239); // @[FFT.scala 34:12]
  wire [31:0] _GEN_241 = 11'hf0 == cnt[10:0] ? $signed(32'sheed9) : $signed(_GEN_240); // @[FFT.scala 34:12]
  wire [31:0] _GEN_242 = 11'hf1 == cnt[10:0] ? $signed(32'sheeb4) : $signed(_GEN_241); // @[FFT.scala 34:12]
  wire [31:0] _GEN_243 = 11'hf2 == cnt[10:0] ? $signed(32'shee90) : $signed(_GEN_242); // @[FFT.scala 34:12]
  wire [31:0] _GEN_244 = 11'hf3 == cnt[10:0] ? $signed(32'shee6b) : $signed(_GEN_243); // @[FFT.scala 34:12]
  wire [31:0] _GEN_245 = 11'hf4 == cnt[10:0] ? $signed(32'shee47) : $signed(_GEN_244); // @[FFT.scala 34:12]
  wire [31:0] _GEN_246 = 11'hf5 == cnt[10:0] ? $signed(32'shee22) : $signed(_GEN_245); // @[FFT.scala 34:12]
  wire [31:0] _GEN_247 = 11'hf6 == cnt[10:0] ? $signed(32'shedfd) : $signed(_GEN_246); // @[FFT.scala 34:12]
  wire [31:0] _GEN_248 = 11'hf7 == cnt[10:0] ? $signed(32'shedd8) : $signed(_GEN_247); // @[FFT.scala 34:12]
  wire [31:0] _GEN_249 = 11'hf8 == cnt[10:0] ? $signed(32'shedb3) : $signed(_GEN_248); // @[FFT.scala 34:12]
  wire [31:0] _GEN_250 = 11'hf9 == cnt[10:0] ? $signed(32'shed8d) : $signed(_GEN_249); // @[FFT.scala 34:12]
  wire [31:0] _GEN_251 = 11'hfa == cnt[10:0] ? $signed(32'shed68) : $signed(_GEN_250); // @[FFT.scala 34:12]
  wire [31:0] _GEN_252 = 11'hfb == cnt[10:0] ? $signed(32'shed42) : $signed(_GEN_251); // @[FFT.scala 34:12]
  wire [31:0] _GEN_253 = 11'hfc == cnt[10:0] ? $signed(32'shed1c) : $signed(_GEN_252); // @[FFT.scala 34:12]
  wire [31:0] _GEN_254 = 11'hfd == cnt[10:0] ? $signed(32'shecf6) : $signed(_GEN_253); // @[FFT.scala 34:12]
  wire [31:0] _GEN_255 = 11'hfe == cnt[10:0] ? $signed(32'shecd0) : $signed(_GEN_254); // @[FFT.scala 34:12]
  wire [31:0] _GEN_256 = 11'hff == cnt[10:0] ? $signed(32'shecaa) : $signed(_GEN_255); // @[FFT.scala 34:12]
  wire [31:0] _GEN_257 = 11'h100 == cnt[10:0] ? $signed(32'shec83) : $signed(_GEN_256); // @[FFT.scala 34:12]
  wire [31:0] _GEN_258 = 11'h101 == cnt[10:0] ? $signed(32'shec5d) : $signed(_GEN_257); // @[FFT.scala 34:12]
  wire [31:0] _GEN_259 = 11'h102 == cnt[10:0] ? $signed(32'shec36) : $signed(_GEN_258); // @[FFT.scala 34:12]
  wire [31:0] _GEN_260 = 11'h103 == cnt[10:0] ? $signed(32'shec0f) : $signed(_GEN_259); // @[FFT.scala 34:12]
  wire [31:0] _GEN_261 = 11'h104 == cnt[10:0] ? $signed(32'shebe8) : $signed(_GEN_260); // @[FFT.scala 34:12]
  wire [31:0] _GEN_262 = 11'h105 == cnt[10:0] ? $signed(32'shebc1) : $signed(_GEN_261); // @[FFT.scala 34:12]
  wire [31:0] _GEN_263 = 11'h106 == cnt[10:0] ? $signed(32'sheb9a) : $signed(_GEN_262); // @[FFT.scala 34:12]
  wire [31:0] _GEN_264 = 11'h107 == cnt[10:0] ? $signed(32'sheb73) : $signed(_GEN_263); // @[FFT.scala 34:12]
  wire [31:0] _GEN_265 = 11'h108 == cnt[10:0] ? $signed(32'sheb4b) : $signed(_GEN_264); // @[FFT.scala 34:12]
  wire [31:0] _GEN_266 = 11'h109 == cnt[10:0] ? $signed(32'sheb23) : $signed(_GEN_265); // @[FFT.scala 34:12]
  wire [31:0] _GEN_267 = 11'h10a == cnt[10:0] ? $signed(32'sheafc) : $signed(_GEN_266); // @[FFT.scala 34:12]
  wire [31:0] _GEN_268 = 11'h10b == cnt[10:0] ? $signed(32'shead4) : $signed(_GEN_267); // @[FFT.scala 34:12]
  wire [31:0] _GEN_269 = 11'h10c == cnt[10:0] ? $signed(32'sheaab) : $signed(_GEN_268); // @[FFT.scala 34:12]
  wire [31:0] _GEN_270 = 11'h10d == cnt[10:0] ? $signed(32'shea83) : $signed(_GEN_269); // @[FFT.scala 34:12]
  wire [31:0] _GEN_271 = 11'h10e == cnt[10:0] ? $signed(32'shea5b) : $signed(_GEN_270); // @[FFT.scala 34:12]
  wire [31:0] _GEN_272 = 11'h10f == cnt[10:0] ? $signed(32'shea32) : $signed(_GEN_271); // @[FFT.scala 34:12]
  wire [31:0] _GEN_273 = 11'h110 == cnt[10:0] ? $signed(32'shea0a) : $signed(_GEN_272); // @[FFT.scala 34:12]
  wire [31:0] _GEN_274 = 11'h111 == cnt[10:0] ? $signed(32'she9e1) : $signed(_GEN_273); // @[FFT.scala 34:12]
  wire [31:0] _GEN_275 = 11'h112 == cnt[10:0] ? $signed(32'she9b8) : $signed(_GEN_274); // @[FFT.scala 34:12]
  wire [31:0] _GEN_276 = 11'h113 == cnt[10:0] ? $signed(32'she98f) : $signed(_GEN_275); // @[FFT.scala 34:12]
  wire [31:0] _GEN_277 = 11'h114 == cnt[10:0] ? $signed(32'she966) : $signed(_GEN_276); // @[FFT.scala 34:12]
  wire [31:0] _GEN_278 = 11'h115 == cnt[10:0] ? $signed(32'she93c) : $signed(_GEN_277); // @[FFT.scala 34:12]
  wire [31:0] _GEN_279 = 11'h116 == cnt[10:0] ? $signed(32'she913) : $signed(_GEN_278); // @[FFT.scala 34:12]
  wire [31:0] _GEN_280 = 11'h117 == cnt[10:0] ? $signed(32'she8e9) : $signed(_GEN_279); // @[FFT.scala 34:12]
  wire [31:0] _GEN_281 = 11'h118 == cnt[10:0] ? $signed(32'she8bf) : $signed(_GEN_280); // @[FFT.scala 34:12]
  wire [31:0] _GEN_282 = 11'h119 == cnt[10:0] ? $signed(32'she895) : $signed(_GEN_281); // @[FFT.scala 34:12]
  wire [31:0] _GEN_283 = 11'h11a == cnt[10:0] ? $signed(32'she86b) : $signed(_GEN_282); // @[FFT.scala 34:12]
  wire [31:0] _GEN_284 = 11'h11b == cnt[10:0] ? $signed(32'she841) : $signed(_GEN_283); // @[FFT.scala 34:12]
  wire [31:0] _GEN_285 = 11'h11c == cnt[10:0] ? $signed(32'she817) : $signed(_GEN_284); // @[FFT.scala 34:12]
  wire [31:0] _GEN_286 = 11'h11d == cnt[10:0] ? $signed(32'she7ec) : $signed(_GEN_285); // @[FFT.scala 34:12]
  wire [31:0] _GEN_287 = 11'h11e == cnt[10:0] ? $signed(32'she7c2) : $signed(_GEN_286); // @[FFT.scala 34:12]
  wire [31:0] _GEN_288 = 11'h11f == cnt[10:0] ? $signed(32'she797) : $signed(_GEN_287); // @[FFT.scala 34:12]
  wire [31:0] _GEN_289 = 11'h120 == cnt[10:0] ? $signed(32'she76c) : $signed(_GEN_288); // @[FFT.scala 34:12]
  wire [31:0] _GEN_290 = 11'h121 == cnt[10:0] ? $signed(32'she741) : $signed(_GEN_289); // @[FFT.scala 34:12]
  wire [31:0] _GEN_291 = 11'h122 == cnt[10:0] ? $signed(32'she716) : $signed(_GEN_290); // @[FFT.scala 34:12]
  wire [31:0] _GEN_292 = 11'h123 == cnt[10:0] ? $signed(32'she6ea) : $signed(_GEN_291); // @[FFT.scala 34:12]
  wire [31:0] _GEN_293 = 11'h124 == cnt[10:0] ? $signed(32'she6bf) : $signed(_GEN_292); // @[FFT.scala 34:12]
  wire [31:0] _GEN_294 = 11'h125 == cnt[10:0] ? $signed(32'she693) : $signed(_GEN_293); // @[FFT.scala 34:12]
  wire [31:0] _GEN_295 = 11'h126 == cnt[10:0] ? $signed(32'she667) : $signed(_GEN_294); // @[FFT.scala 34:12]
  wire [31:0] _GEN_296 = 11'h127 == cnt[10:0] ? $signed(32'she63c) : $signed(_GEN_295); // @[FFT.scala 34:12]
  wire [31:0] _GEN_297 = 11'h128 == cnt[10:0] ? $signed(32'she610) : $signed(_GEN_296); // @[FFT.scala 34:12]
  wire [31:0] _GEN_298 = 11'h129 == cnt[10:0] ? $signed(32'she5e3) : $signed(_GEN_297); // @[FFT.scala 34:12]
  wire [31:0] _GEN_299 = 11'h12a == cnt[10:0] ? $signed(32'she5b7) : $signed(_GEN_298); // @[FFT.scala 34:12]
  wire [31:0] _GEN_300 = 11'h12b == cnt[10:0] ? $signed(32'she58b) : $signed(_GEN_299); // @[FFT.scala 34:12]
  wire [31:0] _GEN_301 = 11'h12c == cnt[10:0] ? $signed(32'she55e) : $signed(_GEN_300); // @[FFT.scala 34:12]
  wire [31:0] _GEN_302 = 11'h12d == cnt[10:0] ? $signed(32'she531) : $signed(_GEN_301); // @[FFT.scala 34:12]
  wire [31:0] _GEN_303 = 11'h12e == cnt[10:0] ? $signed(32'she504) : $signed(_GEN_302); // @[FFT.scala 34:12]
  wire [31:0] _GEN_304 = 11'h12f == cnt[10:0] ? $signed(32'she4d7) : $signed(_GEN_303); // @[FFT.scala 34:12]
  wire [31:0] _GEN_305 = 11'h130 == cnt[10:0] ? $signed(32'she4aa) : $signed(_GEN_304); // @[FFT.scala 34:12]
  wire [31:0] _GEN_306 = 11'h131 == cnt[10:0] ? $signed(32'she47d) : $signed(_GEN_305); // @[FFT.scala 34:12]
  wire [31:0] _GEN_307 = 11'h132 == cnt[10:0] ? $signed(32'she450) : $signed(_GEN_306); // @[FFT.scala 34:12]
  wire [31:0] _GEN_308 = 11'h133 == cnt[10:0] ? $signed(32'she422) : $signed(_GEN_307); // @[FFT.scala 34:12]
  wire [31:0] _GEN_309 = 11'h134 == cnt[10:0] ? $signed(32'she3f4) : $signed(_GEN_308); // @[FFT.scala 34:12]
  wire [31:0] _GEN_310 = 11'h135 == cnt[10:0] ? $signed(32'she3c7) : $signed(_GEN_309); // @[FFT.scala 34:12]
  wire [31:0] _GEN_311 = 11'h136 == cnt[10:0] ? $signed(32'she399) : $signed(_GEN_310); // @[FFT.scala 34:12]
  wire [31:0] _GEN_312 = 11'h137 == cnt[10:0] ? $signed(32'she36b) : $signed(_GEN_311); // @[FFT.scala 34:12]
  wire [31:0] _GEN_313 = 11'h138 == cnt[10:0] ? $signed(32'she33c) : $signed(_GEN_312); // @[FFT.scala 34:12]
  wire [31:0] _GEN_314 = 11'h139 == cnt[10:0] ? $signed(32'she30e) : $signed(_GEN_313); // @[FFT.scala 34:12]
  wire [31:0] _GEN_315 = 11'h13a == cnt[10:0] ? $signed(32'she2df) : $signed(_GEN_314); // @[FFT.scala 34:12]
  wire [31:0] _GEN_316 = 11'h13b == cnt[10:0] ? $signed(32'she2b1) : $signed(_GEN_315); // @[FFT.scala 34:12]
  wire [31:0] _GEN_317 = 11'h13c == cnt[10:0] ? $signed(32'she282) : $signed(_GEN_316); // @[FFT.scala 34:12]
  wire [31:0] _GEN_318 = 11'h13d == cnt[10:0] ? $signed(32'she253) : $signed(_GEN_317); // @[FFT.scala 34:12]
  wire [31:0] _GEN_319 = 11'h13e == cnt[10:0] ? $signed(32'she224) : $signed(_GEN_318); // @[FFT.scala 34:12]
  wire [31:0] _GEN_320 = 11'h13f == cnt[10:0] ? $signed(32'she1f5) : $signed(_GEN_319); // @[FFT.scala 34:12]
  wire [31:0] _GEN_321 = 11'h140 == cnt[10:0] ? $signed(32'she1c6) : $signed(_GEN_320); // @[FFT.scala 34:12]
  wire [31:0] _GEN_322 = 11'h141 == cnt[10:0] ? $signed(32'she196) : $signed(_GEN_321); // @[FFT.scala 34:12]
  wire [31:0] _GEN_323 = 11'h142 == cnt[10:0] ? $signed(32'she167) : $signed(_GEN_322); // @[FFT.scala 34:12]
  wire [31:0] _GEN_324 = 11'h143 == cnt[10:0] ? $signed(32'she137) : $signed(_GEN_323); // @[FFT.scala 34:12]
  wire [31:0] _GEN_325 = 11'h144 == cnt[10:0] ? $signed(32'she107) : $signed(_GEN_324); // @[FFT.scala 34:12]
  wire [31:0] _GEN_326 = 11'h145 == cnt[10:0] ? $signed(32'she0d7) : $signed(_GEN_325); // @[FFT.scala 34:12]
  wire [31:0] _GEN_327 = 11'h146 == cnt[10:0] ? $signed(32'she0a7) : $signed(_GEN_326); // @[FFT.scala 34:12]
  wire [31:0] _GEN_328 = 11'h147 == cnt[10:0] ? $signed(32'she077) : $signed(_GEN_327); // @[FFT.scala 34:12]
  wire [31:0] _GEN_329 = 11'h148 == cnt[10:0] ? $signed(32'she046) : $signed(_GEN_328); // @[FFT.scala 34:12]
  wire [31:0] _GEN_330 = 11'h149 == cnt[10:0] ? $signed(32'she016) : $signed(_GEN_329); // @[FFT.scala 34:12]
  wire [31:0] _GEN_331 = 11'h14a == cnt[10:0] ? $signed(32'shdfe5) : $signed(_GEN_330); // @[FFT.scala 34:12]
  wire [31:0] _GEN_332 = 11'h14b == cnt[10:0] ? $signed(32'shdfb4) : $signed(_GEN_331); // @[FFT.scala 34:12]
  wire [31:0] _GEN_333 = 11'h14c == cnt[10:0] ? $signed(32'shdf83) : $signed(_GEN_332); // @[FFT.scala 34:12]
  wire [31:0] _GEN_334 = 11'h14d == cnt[10:0] ? $signed(32'shdf52) : $signed(_GEN_333); // @[FFT.scala 34:12]
  wire [31:0] _GEN_335 = 11'h14e == cnt[10:0] ? $signed(32'shdf21) : $signed(_GEN_334); // @[FFT.scala 34:12]
  wire [31:0] _GEN_336 = 11'h14f == cnt[10:0] ? $signed(32'shdef0) : $signed(_GEN_335); // @[FFT.scala 34:12]
  wire [31:0] _GEN_337 = 11'h150 == cnt[10:0] ? $signed(32'shdebe) : $signed(_GEN_336); // @[FFT.scala 34:12]
  wire [31:0] _GEN_338 = 11'h151 == cnt[10:0] ? $signed(32'shde8c) : $signed(_GEN_337); // @[FFT.scala 34:12]
  wire [31:0] _GEN_339 = 11'h152 == cnt[10:0] ? $signed(32'shde5b) : $signed(_GEN_338); // @[FFT.scala 34:12]
  wire [31:0] _GEN_340 = 11'h153 == cnt[10:0] ? $signed(32'shde29) : $signed(_GEN_339); // @[FFT.scala 34:12]
  wire [31:0] _GEN_341 = 11'h154 == cnt[10:0] ? $signed(32'shddf7) : $signed(_GEN_340); // @[FFT.scala 34:12]
  wire [31:0] _GEN_342 = 11'h155 == cnt[10:0] ? $signed(32'shddc5) : $signed(_GEN_341); // @[FFT.scala 34:12]
  wire [31:0] _GEN_343 = 11'h156 == cnt[10:0] ? $signed(32'shdd92) : $signed(_GEN_342); // @[FFT.scala 34:12]
  wire [31:0] _GEN_344 = 11'h157 == cnt[10:0] ? $signed(32'shdd60) : $signed(_GEN_343); // @[FFT.scala 34:12]
  wire [31:0] _GEN_345 = 11'h158 == cnt[10:0] ? $signed(32'shdd2d) : $signed(_GEN_344); // @[FFT.scala 34:12]
  wire [31:0] _GEN_346 = 11'h159 == cnt[10:0] ? $signed(32'shdcfb) : $signed(_GEN_345); // @[FFT.scala 34:12]
  wire [31:0] _GEN_347 = 11'h15a == cnt[10:0] ? $signed(32'shdcc8) : $signed(_GEN_346); // @[FFT.scala 34:12]
  wire [31:0] _GEN_348 = 11'h15b == cnt[10:0] ? $signed(32'shdc95) : $signed(_GEN_347); // @[FFT.scala 34:12]
  wire [31:0] _GEN_349 = 11'h15c == cnt[10:0] ? $signed(32'shdc62) : $signed(_GEN_348); // @[FFT.scala 34:12]
  wire [31:0] _GEN_350 = 11'h15d == cnt[10:0] ? $signed(32'shdc2f) : $signed(_GEN_349); // @[FFT.scala 34:12]
  wire [31:0] _GEN_351 = 11'h15e == cnt[10:0] ? $signed(32'shdbfb) : $signed(_GEN_350); // @[FFT.scala 34:12]
  wire [31:0] _GEN_352 = 11'h15f == cnt[10:0] ? $signed(32'shdbc8) : $signed(_GEN_351); // @[FFT.scala 34:12]
  wire [31:0] _GEN_353 = 11'h160 == cnt[10:0] ? $signed(32'shdb94) : $signed(_GEN_352); // @[FFT.scala 34:12]
  wire [31:0] _GEN_354 = 11'h161 == cnt[10:0] ? $signed(32'shdb60) : $signed(_GEN_353); // @[FFT.scala 34:12]
  wire [31:0] _GEN_355 = 11'h162 == cnt[10:0] ? $signed(32'shdb2c) : $signed(_GEN_354); // @[FFT.scala 34:12]
  wire [31:0] _GEN_356 = 11'h163 == cnt[10:0] ? $signed(32'shdaf8) : $signed(_GEN_355); // @[FFT.scala 34:12]
  wire [31:0] _GEN_357 = 11'h164 == cnt[10:0] ? $signed(32'shdac4) : $signed(_GEN_356); // @[FFT.scala 34:12]
  wire [31:0] _GEN_358 = 11'h165 == cnt[10:0] ? $signed(32'shda90) : $signed(_GEN_357); // @[FFT.scala 34:12]
  wire [31:0] _GEN_359 = 11'h166 == cnt[10:0] ? $signed(32'shda5c) : $signed(_GEN_358); // @[FFT.scala 34:12]
  wire [31:0] _GEN_360 = 11'h167 == cnt[10:0] ? $signed(32'shda27) : $signed(_GEN_359); // @[FFT.scala 34:12]
  wire [31:0] _GEN_361 = 11'h168 == cnt[10:0] ? $signed(32'shd9f2) : $signed(_GEN_360); // @[FFT.scala 34:12]
  wire [31:0] _GEN_362 = 11'h169 == cnt[10:0] ? $signed(32'shd9be) : $signed(_GEN_361); // @[FFT.scala 34:12]
  wire [31:0] _GEN_363 = 11'h16a == cnt[10:0] ? $signed(32'shd989) : $signed(_GEN_362); // @[FFT.scala 34:12]
  wire [31:0] _GEN_364 = 11'h16b == cnt[10:0] ? $signed(32'shd954) : $signed(_GEN_363); // @[FFT.scala 34:12]
  wire [31:0] _GEN_365 = 11'h16c == cnt[10:0] ? $signed(32'shd91e) : $signed(_GEN_364); // @[FFT.scala 34:12]
  wire [31:0] _GEN_366 = 11'h16d == cnt[10:0] ? $signed(32'shd8e9) : $signed(_GEN_365); // @[FFT.scala 34:12]
  wire [31:0] _GEN_367 = 11'h16e == cnt[10:0] ? $signed(32'shd8b4) : $signed(_GEN_366); // @[FFT.scala 34:12]
  wire [31:0] _GEN_368 = 11'h16f == cnt[10:0] ? $signed(32'shd87e) : $signed(_GEN_367); // @[FFT.scala 34:12]
  wire [31:0] _GEN_369 = 11'h170 == cnt[10:0] ? $signed(32'shd848) : $signed(_GEN_368); // @[FFT.scala 34:12]
  wire [31:0] _GEN_370 = 11'h171 == cnt[10:0] ? $signed(32'shd812) : $signed(_GEN_369); // @[FFT.scala 34:12]
  wire [31:0] _GEN_371 = 11'h172 == cnt[10:0] ? $signed(32'shd7dc) : $signed(_GEN_370); // @[FFT.scala 34:12]
  wire [31:0] _GEN_372 = 11'h173 == cnt[10:0] ? $signed(32'shd7a6) : $signed(_GEN_371); // @[FFT.scala 34:12]
  wire [31:0] _GEN_373 = 11'h174 == cnt[10:0] ? $signed(32'shd770) : $signed(_GEN_372); // @[FFT.scala 34:12]
  wire [31:0] _GEN_374 = 11'h175 == cnt[10:0] ? $signed(32'shd73a) : $signed(_GEN_373); // @[FFT.scala 34:12]
  wire [31:0] _GEN_375 = 11'h176 == cnt[10:0] ? $signed(32'shd703) : $signed(_GEN_374); // @[FFT.scala 34:12]
  wire [31:0] _GEN_376 = 11'h177 == cnt[10:0] ? $signed(32'shd6cd) : $signed(_GEN_375); // @[FFT.scala 34:12]
  wire [31:0] _GEN_377 = 11'h178 == cnt[10:0] ? $signed(32'shd696) : $signed(_GEN_376); // @[FFT.scala 34:12]
  wire [31:0] _GEN_378 = 11'h179 == cnt[10:0] ? $signed(32'shd65f) : $signed(_GEN_377); // @[FFT.scala 34:12]
  wire [31:0] _GEN_379 = 11'h17a == cnt[10:0] ? $signed(32'shd628) : $signed(_GEN_378); // @[FFT.scala 34:12]
  wire [31:0] _GEN_380 = 11'h17b == cnt[10:0] ? $signed(32'shd5f1) : $signed(_GEN_379); // @[FFT.scala 34:12]
  wire [31:0] _GEN_381 = 11'h17c == cnt[10:0] ? $signed(32'shd5ba) : $signed(_GEN_380); // @[FFT.scala 34:12]
  wire [31:0] _GEN_382 = 11'h17d == cnt[10:0] ? $signed(32'shd582) : $signed(_GEN_381); // @[FFT.scala 34:12]
  wire [31:0] _GEN_383 = 11'h17e == cnt[10:0] ? $signed(32'shd54b) : $signed(_GEN_382); // @[FFT.scala 34:12]
  wire [31:0] _GEN_384 = 11'h17f == cnt[10:0] ? $signed(32'shd513) : $signed(_GEN_383); // @[FFT.scala 34:12]
  wire [31:0] _GEN_385 = 11'h180 == cnt[10:0] ? $signed(32'shd4db) : $signed(_GEN_384); // @[FFT.scala 34:12]
  wire [31:0] _GEN_386 = 11'h181 == cnt[10:0] ? $signed(32'shd4a3) : $signed(_GEN_385); // @[FFT.scala 34:12]
  wire [31:0] _GEN_387 = 11'h182 == cnt[10:0] ? $signed(32'shd46b) : $signed(_GEN_386); // @[FFT.scala 34:12]
  wire [31:0] _GEN_388 = 11'h183 == cnt[10:0] ? $signed(32'shd433) : $signed(_GEN_387); // @[FFT.scala 34:12]
  wire [31:0] _GEN_389 = 11'h184 == cnt[10:0] ? $signed(32'shd3fb) : $signed(_GEN_388); // @[FFT.scala 34:12]
  wire [31:0] _GEN_390 = 11'h185 == cnt[10:0] ? $signed(32'shd3c2) : $signed(_GEN_389); // @[FFT.scala 34:12]
  wire [31:0] _GEN_391 = 11'h186 == cnt[10:0] ? $signed(32'shd38a) : $signed(_GEN_390); // @[FFT.scala 34:12]
  wire [31:0] _GEN_392 = 11'h187 == cnt[10:0] ? $signed(32'shd351) : $signed(_GEN_391); // @[FFT.scala 34:12]
  wire [31:0] _GEN_393 = 11'h188 == cnt[10:0] ? $signed(32'shd318) : $signed(_GEN_392); // @[FFT.scala 34:12]
  wire [31:0] _GEN_394 = 11'h189 == cnt[10:0] ? $signed(32'shd2df) : $signed(_GEN_393); // @[FFT.scala 34:12]
  wire [31:0] _GEN_395 = 11'h18a == cnt[10:0] ? $signed(32'shd2a6) : $signed(_GEN_394); // @[FFT.scala 34:12]
  wire [31:0] _GEN_396 = 11'h18b == cnt[10:0] ? $signed(32'shd26d) : $signed(_GEN_395); // @[FFT.scala 34:12]
  wire [31:0] _GEN_397 = 11'h18c == cnt[10:0] ? $signed(32'shd234) : $signed(_GEN_396); // @[FFT.scala 34:12]
  wire [31:0] _GEN_398 = 11'h18d == cnt[10:0] ? $signed(32'shd1fa) : $signed(_GEN_397); // @[FFT.scala 34:12]
  wire [31:0] _GEN_399 = 11'h18e == cnt[10:0] ? $signed(32'shd1c1) : $signed(_GEN_398); // @[FFT.scala 34:12]
  wire [31:0] _GEN_400 = 11'h18f == cnt[10:0] ? $signed(32'shd187) : $signed(_GEN_399); // @[FFT.scala 34:12]
  wire [31:0] _GEN_401 = 11'h190 == cnt[10:0] ? $signed(32'shd14d) : $signed(_GEN_400); // @[FFT.scala 34:12]
  wire [31:0] _GEN_402 = 11'h191 == cnt[10:0] ? $signed(32'shd113) : $signed(_GEN_401); // @[FFT.scala 34:12]
  wire [31:0] _GEN_403 = 11'h192 == cnt[10:0] ? $signed(32'shd0d9) : $signed(_GEN_402); // @[FFT.scala 34:12]
  wire [31:0] _GEN_404 = 11'h193 == cnt[10:0] ? $signed(32'shd09f) : $signed(_GEN_403); // @[FFT.scala 34:12]
  wire [31:0] _GEN_405 = 11'h194 == cnt[10:0] ? $signed(32'shd065) : $signed(_GEN_404); // @[FFT.scala 34:12]
  wire [31:0] _GEN_406 = 11'h195 == cnt[10:0] ? $signed(32'shd02a) : $signed(_GEN_405); // @[FFT.scala 34:12]
  wire [31:0] _GEN_407 = 11'h196 == cnt[10:0] ? $signed(32'shcff0) : $signed(_GEN_406); // @[FFT.scala 34:12]
  wire [31:0] _GEN_408 = 11'h197 == cnt[10:0] ? $signed(32'shcfb5) : $signed(_GEN_407); // @[FFT.scala 34:12]
  wire [31:0] _GEN_409 = 11'h198 == cnt[10:0] ? $signed(32'shcf7a) : $signed(_GEN_408); // @[FFT.scala 34:12]
  wire [31:0] _GEN_410 = 11'h199 == cnt[10:0] ? $signed(32'shcf3f) : $signed(_GEN_409); // @[FFT.scala 34:12]
  wire [31:0] _GEN_411 = 11'h19a == cnt[10:0] ? $signed(32'shcf04) : $signed(_GEN_410); // @[FFT.scala 34:12]
  wire [31:0] _GEN_412 = 11'h19b == cnt[10:0] ? $signed(32'shcec9) : $signed(_GEN_411); // @[FFT.scala 34:12]
  wire [31:0] _GEN_413 = 11'h19c == cnt[10:0] ? $signed(32'shce8e) : $signed(_GEN_412); // @[FFT.scala 34:12]
  wire [31:0] _GEN_414 = 11'h19d == cnt[10:0] ? $signed(32'shce52) : $signed(_GEN_413); // @[FFT.scala 34:12]
  wire [31:0] _GEN_415 = 11'h19e == cnt[10:0] ? $signed(32'shce17) : $signed(_GEN_414); // @[FFT.scala 34:12]
  wire [31:0] _GEN_416 = 11'h19f == cnt[10:0] ? $signed(32'shcddb) : $signed(_GEN_415); // @[FFT.scala 34:12]
  wire [31:0] _GEN_417 = 11'h1a0 == cnt[10:0] ? $signed(32'shcd9f) : $signed(_GEN_416); // @[FFT.scala 34:12]
  wire [31:0] _GEN_418 = 11'h1a1 == cnt[10:0] ? $signed(32'shcd63) : $signed(_GEN_417); // @[FFT.scala 34:12]
  wire [31:0] _GEN_419 = 11'h1a2 == cnt[10:0] ? $signed(32'shcd27) : $signed(_GEN_418); // @[FFT.scala 34:12]
  wire [31:0] _GEN_420 = 11'h1a3 == cnt[10:0] ? $signed(32'shcceb) : $signed(_GEN_419); // @[FFT.scala 34:12]
  wire [31:0] _GEN_421 = 11'h1a4 == cnt[10:0] ? $signed(32'shccae) : $signed(_GEN_420); // @[FFT.scala 34:12]
  wire [31:0] _GEN_422 = 11'h1a5 == cnt[10:0] ? $signed(32'shcc72) : $signed(_GEN_421); // @[FFT.scala 34:12]
  wire [31:0] _GEN_423 = 11'h1a6 == cnt[10:0] ? $signed(32'shcc35) : $signed(_GEN_422); // @[FFT.scala 34:12]
  wire [31:0] _GEN_424 = 11'h1a7 == cnt[10:0] ? $signed(32'shcbf9) : $signed(_GEN_423); // @[FFT.scala 34:12]
  wire [31:0] _GEN_425 = 11'h1a8 == cnt[10:0] ? $signed(32'shcbbc) : $signed(_GEN_424); // @[FFT.scala 34:12]
  wire [31:0] _GEN_426 = 11'h1a9 == cnt[10:0] ? $signed(32'shcb7f) : $signed(_GEN_425); // @[FFT.scala 34:12]
  wire [31:0] _GEN_427 = 11'h1aa == cnt[10:0] ? $signed(32'shcb42) : $signed(_GEN_426); // @[FFT.scala 34:12]
  wire [31:0] _GEN_428 = 11'h1ab == cnt[10:0] ? $signed(32'shcb05) : $signed(_GEN_427); // @[FFT.scala 34:12]
  wire [31:0] _GEN_429 = 11'h1ac == cnt[10:0] ? $signed(32'shcac7) : $signed(_GEN_428); // @[FFT.scala 34:12]
  wire [31:0] _GEN_430 = 11'h1ad == cnt[10:0] ? $signed(32'shca8a) : $signed(_GEN_429); // @[FFT.scala 34:12]
  wire [31:0] _GEN_431 = 11'h1ae == cnt[10:0] ? $signed(32'shca4d) : $signed(_GEN_430); // @[FFT.scala 34:12]
  wire [31:0] _GEN_432 = 11'h1af == cnt[10:0] ? $signed(32'shca0f) : $signed(_GEN_431); // @[FFT.scala 34:12]
  wire [31:0] _GEN_433 = 11'h1b0 == cnt[10:0] ? $signed(32'shc9d1) : $signed(_GEN_432); // @[FFT.scala 34:12]
  wire [31:0] _GEN_434 = 11'h1b1 == cnt[10:0] ? $signed(32'shc993) : $signed(_GEN_433); // @[FFT.scala 34:12]
  wire [31:0] _GEN_435 = 11'h1b2 == cnt[10:0] ? $signed(32'shc955) : $signed(_GEN_434); // @[FFT.scala 34:12]
  wire [31:0] _GEN_436 = 11'h1b3 == cnt[10:0] ? $signed(32'shc917) : $signed(_GEN_435); // @[FFT.scala 34:12]
  wire [31:0] _GEN_437 = 11'h1b4 == cnt[10:0] ? $signed(32'shc8d9) : $signed(_GEN_436); // @[FFT.scala 34:12]
  wire [31:0] _GEN_438 = 11'h1b5 == cnt[10:0] ? $signed(32'shc89a) : $signed(_GEN_437); // @[FFT.scala 34:12]
  wire [31:0] _GEN_439 = 11'h1b6 == cnt[10:0] ? $signed(32'shc85c) : $signed(_GEN_438); // @[FFT.scala 34:12]
  wire [31:0] _GEN_440 = 11'h1b7 == cnt[10:0] ? $signed(32'shc81d) : $signed(_GEN_439); // @[FFT.scala 34:12]
  wire [31:0] _GEN_441 = 11'h1b8 == cnt[10:0] ? $signed(32'shc7de) : $signed(_GEN_440); // @[FFT.scala 34:12]
  wire [31:0] _GEN_442 = 11'h1b9 == cnt[10:0] ? $signed(32'shc7a0) : $signed(_GEN_441); // @[FFT.scala 34:12]
  wire [31:0] _GEN_443 = 11'h1ba == cnt[10:0] ? $signed(32'shc761) : $signed(_GEN_442); // @[FFT.scala 34:12]
  wire [31:0] _GEN_444 = 11'h1bb == cnt[10:0] ? $signed(32'shc721) : $signed(_GEN_443); // @[FFT.scala 34:12]
  wire [31:0] _GEN_445 = 11'h1bc == cnt[10:0] ? $signed(32'shc6e2) : $signed(_GEN_444); // @[FFT.scala 34:12]
  wire [31:0] _GEN_446 = 11'h1bd == cnt[10:0] ? $signed(32'shc6a3) : $signed(_GEN_445); // @[FFT.scala 34:12]
  wire [31:0] _GEN_447 = 11'h1be == cnt[10:0] ? $signed(32'shc663) : $signed(_GEN_446); // @[FFT.scala 34:12]
  wire [31:0] _GEN_448 = 11'h1bf == cnt[10:0] ? $signed(32'shc624) : $signed(_GEN_447); // @[FFT.scala 34:12]
  wire [31:0] _GEN_449 = 11'h1c0 == cnt[10:0] ? $signed(32'shc5e4) : $signed(_GEN_448); // @[FFT.scala 34:12]
  wire [31:0] _GEN_450 = 11'h1c1 == cnt[10:0] ? $signed(32'shc5a4) : $signed(_GEN_449); // @[FFT.scala 34:12]
  wire [31:0] _GEN_451 = 11'h1c2 == cnt[10:0] ? $signed(32'shc564) : $signed(_GEN_450); // @[FFT.scala 34:12]
  wire [31:0] _GEN_452 = 11'h1c3 == cnt[10:0] ? $signed(32'shc524) : $signed(_GEN_451); // @[FFT.scala 34:12]
  wire [31:0] _GEN_453 = 11'h1c4 == cnt[10:0] ? $signed(32'shc4e4) : $signed(_GEN_452); // @[FFT.scala 34:12]
  wire [31:0] _GEN_454 = 11'h1c5 == cnt[10:0] ? $signed(32'shc4a4) : $signed(_GEN_453); // @[FFT.scala 34:12]
  wire [31:0] _GEN_455 = 11'h1c6 == cnt[10:0] ? $signed(32'shc463) : $signed(_GEN_454); // @[FFT.scala 34:12]
  wire [31:0] _GEN_456 = 11'h1c7 == cnt[10:0] ? $signed(32'shc423) : $signed(_GEN_455); // @[FFT.scala 34:12]
  wire [31:0] _GEN_457 = 11'h1c8 == cnt[10:0] ? $signed(32'shc3e2) : $signed(_GEN_456); // @[FFT.scala 34:12]
  wire [31:0] _GEN_458 = 11'h1c9 == cnt[10:0] ? $signed(32'shc3a1) : $signed(_GEN_457); // @[FFT.scala 34:12]
  wire [31:0] _GEN_459 = 11'h1ca == cnt[10:0] ? $signed(32'shc360) : $signed(_GEN_458); // @[FFT.scala 34:12]
  wire [31:0] _GEN_460 = 11'h1cb == cnt[10:0] ? $signed(32'shc31f) : $signed(_GEN_459); // @[FFT.scala 34:12]
  wire [31:0] _GEN_461 = 11'h1cc == cnt[10:0] ? $signed(32'shc2de) : $signed(_GEN_460); // @[FFT.scala 34:12]
  wire [31:0] _GEN_462 = 11'h1cd == cnt[10:0] ? $signed(32'shc29d) : $signed(_GEN_461); // @[FFT.scala 34:12]
  wire [31:0] _GEN_463 = 11'h1ce == cnt[10:0] ? $signed(32'shc25c) : $signed(_GEN_462); // @[FFT.scala 34:12]
  wire [31:0] _GEN_464 = 11'h1cf == cnt[10:0] ? $signed(32'shc21a) : $signed(_GEN_463); // @[FFT.scala 34:12]
  wire [31:0] _GEN_465 = 11'h1d0 == cnt[10:0] ? $signed(32'shc1d8) : $signed(_GEN_464); // @[FFT.scala 34:12]
  wire [31:0] _GEN_466 = 11'h1d1 == cnt[10:0] ? $signed(32'shc197) : $signed(_GEN_465); // @[FFT.scala 34:12]
  wire [31:0] _GEN_467 = 11'h1d2 == cnt[10:0] ? $signed(32'shc155) : $signed(_GEN_466); // @[FFT.scala 34:12]
  wire [31:0] _GEN_468 = 11'h1d3 == cnt[10:0] ? $signed(32'shc113) : $signed(_GEN_467); // @[FFT.scala 34:12]
  wire [31:0] _GEN_469 = 11'h1d4 == cnt[10:0] ? $signed(32'shc0d1) : $signed(_GEN_468); // @[FFT.scala 34:12]
  wire [31:0] _GEN_470 = 11'h1d5 == cnt[10:0] ? $signed(32'shc08f) : $signed(_GEN_469); // @[FFT.scala 34:12]
  wire [31:0] _GEN_471 = 11'h1d6 == cnt[10:0] ? $signed(32'shc04c) : $signed(_GEN_470); // @[FFT.scala 34:12]
  wire [31:0] _GEN_472 = 11'h1d7 == cnt[10:0] ? $signed(32'shc00a) : $signed(_GEN_471); // @[FFT.scala 34:12]
  wire [31:0] _GEN_473 = 11'h1d8 == cnt[10:0] ? $signed(32'shbfc7) : $signed(_GEN_472); // @[FFT.scala 34:12]
  wire [31:0] _GEN_474 = 11'h1d9 == cnt[10:0] ? $signed(32'shbf85) : $signed(_GEN_473); // @[FFT.scala 34:12]
  wire [31:0] _GEN_475 = 11'h1da == cnt[10:0] ? $signed(32'shbf42) : $signed(_GEN_474); // @[FFT.scala 34:12]
  wire [31:0] _GEN_476 = 11'h1db == cnt[10:0] ? $signed(32'shbeff) : $signed(_GEN_475); // @[FFT.scala 34:12]
  wire [31:0] _GEN_477 = 11'h1dc == cnt[10:0] ? $signed(32'shbebc) : $signed(_GEN_476); // @[FFT.scala 34:12]
  wire [31:0] _GEN_478 = 11'h1dd == cnt[10:0] ? $signed(32'shbe79) : $signed(_GEN_477); // @[FFT.scala 34:12]
  wire [31:0] _GEN_479 = 11'h1de == cnt[10:0] ? $signed(32'shbe36) : $signed(_GEN_478); // @[FFT.scala 34:12]
  wire [31:0] _GEN_480 = 11'h1df == cnt[10:0] ? $signed(32'shbdf2) : $signed(_GEN_479); // @[FFT.scala 34:12]
  wire [31:0] _GEN_481 = 11'h1e0 == cnt[10:0] ? $signed(32'shbdaf) : $signed(_GEN_480); // @[FFT.scala 34:12]
  wire [31:0] _GEN_482 = 11'h1e1 == cnt[10:0] ? $signed(32'shbd6b) : $signed(_GEN_481); // @[FFT.scala 34:12]
  wire [31:0] _GEN_483 = 11'h1e2 == cnt[10:0] ? $signed(32'shbd28) : $signed(_GEN_482); // @[FFT.scala 34:12]
  wire [31:0] _GEN_484 = 11'h1e3 == cnt[10:0] ? $signed(32'shbce4) : $signed(_GEN_483); // @[FFT.scala 34:12]
  wire [31:0] _GEN_485 = 11'h1e4 == cnt[10:0] ? $signed(32'shbca0) : $signed(_GEN_484); // @[FFT.scala 34:12]
  wire [31:0] _GEN_486 = 11'h1e5 == cnt[10:0] ? $signed(32'shbc5c) : $signed(_GEN_485); // @[FFT.scala 34:12]
  wire [31:0] _GEN_487 = 11'h1e6 == cnt[10:0] ? $signed(32'shbc18) : $signed(_GEN_486); // @[FFT.scala 34:12]
  wire [31:0] _GEN_488 = 11'h1e7 == cnt[10:0] ? $signed(32'shbbd4) : $signed(_GEN_487); // @[FFT.scala 34:12]
  wire [31:0] _GEN_489 = 11'h1e8 == cnt[10:0] ? $signed(32'shbb8f) : $signed(_GEN_488); // @[FFT.scala 34:12]
  wire [31:0] _GEN_490 = 11'h1e9 == cnt[10:0] ? $signed(32'shbb4b) : $signed(_GEN_489); // @[FFT.scala 34:12]
  wire [31:0] _GEN_491 = 11'h1ea == cnt[10:0] ? $signed(32'shbb06) : $signed(_GEN_490); // @[FFT.scala 34:12]
  wire [31:0] _GEN_492 = 11'h1eb == cnt[10:0] ? $signed(32'shbac1) : $signed(_GEN_491); // @[FFT.scala 34:12]
  wire [31:0] _GEN_493 = 11'h1ec == cnt[10:0] ? $signed(32'shba7d) : $signed(_GEN_492); // @[FFT.scala 34:12]
  wire [31:0] _GEN_494 = 11'h1ed == cnt[10:0] ? $signed(32'shba38) : $signed(_GEN_493); // @[FFT.scala 34:12]
  wire [31:0] _GEN_495 = 11'h1ee == cnt[10:0] ? $signed(32'shb9f3) : $signed(_GEN_494); // @[FFT.scala 34:12]
  wire [31:0] _GEN_496 = 11'h1ef == cnt[10:0] ? $signed(32'shb9ae) : $signed(_GEN_495); // @[FFT.scala 34:12]
  wire [31:0] _GEN_497 = 11'h1f0 == cnt[10:0] ? $signed(32'shb968) : $signed(_GEN_496); // @[FFT.scala 34:12]
  wire [31:0] _GEN_498 = 11'h1f1 == cnt[10:0] ? $signed(32'shb923) : $signed(_GEN_497); // @[FFT.scala 34:12]
  wire [31:0] _GEN_499 = 11'h1f2 == cnt[10:0] ? $signed(32'shb8dd) : $signed(_GEN_498); // @[FFT.scala 34:12]
  wire [31:0] _GEN_500 = 11'h1f3 == cnt[10:0] ? $signed(32'shb898) : $signed(_GEN_499); // @[FFT.scala 34:12]
  wire [31:0] _GEN_501 = 11'h1f4 == cnt[10:0] ? $signed(32'shb852) : $signed(_GEN_500); // @[FFT.scala 34:12]
  wire [31:0] _GEN_502 = 11'h1f5 == cnt[10:0] ? $signed(32'shb80c) : $signed(_GEN_501); // @[FFT.scala 34:12]
  wire [31:0] _GEN_503 = 11'h1f6 == cnt[10:0] ? $signed(32'shb7c6) : $signed(_GEN_502); // @[FFT.scala 34:12]
  wire [31:0] _GEN_504 = 11'h1f7 == cnt[10:0] ? $signed(32'shb780) : $signed(_GEN_503); // @[FFT.scala 34:12]
  wire [31:0] _GEN_505 = 11'h1f8 == cnt[10:0] ? $signed(32'shb73a) : $signed(_GEN_504); // @[FFT.scala 34:12]
  wire [31:0] _GEN_506 = 11'h1f9 == cnt[10:0] ? $signed(32'shb6f4) : $signed(_GEN_505); // @[FFT.scala 34:12]
  wire [31:0] _GEN_507 = 11'h1fa == cnt[10:0] ? $signed(32'shb6ad) : $signed(_GEN_506); // @[FFT.scala 34:12]
  wire [31:0] _GEN_508 = 11'h1fb == cnt[10:0] ? $signed(32'shb667) : $signed(_GEN_507); // @[FFT.scala 34:12]
  wire [31:0] _GEN_509 = 11'h1fc == cnt[10:0] ? $signed(32'shb620) : $signed(_GEN_508); // @[FFT.scala 34:12]
  wire [31:0] _GEN_510 = 11'h1fd == cnt[10:0] ? $signed(32'shb5da) : $signed(_GEN_509); // @[FFT.scala 34:12]
  wire [31:0] _GEN_511 = 11'h1fe == cnt[10:0] ? $signed(32'shb593) : $signed(_GEN_510); // @[FFT.scala 34:12]
  wire [31:0] _GEN_512 = 11'h1ff == cnt[10:0] ? $signed(32'shb54c) : $signed(_GEN_511); // @[FFT.scala 34:12]
  wire [31:0] _GEN_513 = 11'h200 == cnt[10:0] ? $signed(32'shb505) : $signed(_GEN_512); // @[FFT.scala 34:12]
  wire [31:0] _GEN_514 = 11'h201 == cnt[10:0] ? $signed(32'shb4be) : $signed(_GEN_513); // @[FFT.scala 34:12]
  wire [31:0] _GEN_515 = 11'h202 == cnt[10:0] ? $signed(32'shb477) : $signed(_GEN_514); // @[FFT.scala 34:12]
  wire [31:0] _GEN_516 = 11'h203 == cnt[10:0] ? $signed(32'shb42f) : $signed(_GEN_515); // @[FFT.scala 34:12]
  wire [31:0] _GEN_517 = 11'h204 == cnt[10:0] ? $signed(32'shb3e8) : $signed(_GEN_516); // @[FFT.scala 34:12]
  wire [31:0] _GEN_518 = 11'h205 == cnt[10:0] ? $signed(32'shb3a0) : $signed(_GEN_517); // @[FFT.scala 34:12]
  wire [31:0] _GEN_519 = 11'h206 == cnt[10:0] ? $signed(32'shb358) : $signed(_GEN_518); // @[FFT.scala 34:12]
  wire [31:0] _GEN_520 = 11'h207 == cnt[10:0] ? $signed(32'shb311) : $signed(_GEN_519); // @[FFT.scala 34:12]
  wire [31:0] _GEN_521 = 11'h208 == cnt[10:0] ? $signed(32'shb2c9) : $signed(_GEN_520); // @[FFT.scala 34:12]
  wire [31:0] _GEN_522 = 11'h209 == cnt[10:0] ? $signed(32'shb281) : $signed(_GEN_521); // @[FFT.scala 34:12]
  wire [31:0] _GEN_523 = 11'h20a == cnt[10:0] ? $signed(32'shb239) : $signed(_GEN_522); // @[FFT.scala 34:12]
  wire [31:0] _GEN_524 = 11'h20b == cnt[10:0] ? $signed(32'shb1f0) : $signed(_GEN_523); // @[FFT.scala 34:12]
  wire [31:0] _GEN_525 = 11'h20c == cnt[10:0] ? $signed(32'shb1a8) : $signed(_GEN_524); // @[FFT.scala 34:12]
  wire [31:0] _GEN_526 = 11'h20d == cnt[10:0] ? $signed(32'shb160) : $signed(_GEN_525); // @[FFT.scala 34:12]
  wire [31:0] _GEN_527 = 11'h20e == cnt[10:0] ? $signed(32'shb117) : $signed(_GEN_526); // @[FFT.scala 34:12]
  wire [31:0] _GEN_528 = 11'h20f == cnt[10:0] ? $signed(32'shb0ce) : $signed(_GEN_527); // @[FFT.scala 34:12]
  wire [31:0] _GEN_529 = 11'h210 == cnt[10:0] ? $signed(32'shb086) : $signed(_GEN_528); // @[FFT.scala 34:12]
  wire [31:0] _GEN_530 = 11'h211 == cnt[10:0] ? $signed(32'shb03d) : $signed(_GEN_529); // @[FFT.scala 34:12]
  wire [31:0] _GEN_531 = 11'h212 == cnt[10:0] ? $signed(32'shaff4) : $signed(_GEN_530); // @[FFT.scala 34:12]
  wire [31:0] _GEN_532 = 11'h213 == cnt[10:0] ? $signed(32'shafab) : $signed(_GEN_531); // @[FFT.scala 34:12]
  wire [31:0] _GEN_533 = 11'h214 == cnt[10:0] ? $signed(32'shaf62) : $signed(_GEN_532); // @[FFT.scala 34:12]
  wire [31:0] _GEN_534 = 11'h215 == cnt[10:0] ? $signed(32'shaf18) : $signed(_GEN_533); // @[FFT.scala 34:12]
  wire [31:0] _GEN_535 = 11'h216 == cnt[10:0] ? $signed(32'shaecf) : $signed(_GEN_534); // @[FFT.scala 34:12]
  wire [31:0] _GEN_536 = 11'h217 == cnt[10:0] ? $signed(32'shae85) : $signed(_GEN_535); // @[FFT.scala 34:12]
  wire [31:0] _GEN_537 = 11'h218 == cnt[10:0] ? $signed(32'shae3c) : $signed(_GEN_536); // @[FFT.scala 34:12]
  wire [31:0] _GEN_538 = 11'h219 == cnt[10:0] ? $signed(32'shadf2) : $signed(_GEN_537); // @[FFT.scala 34:12]
  wire [31:0] _GEN_539 = 11'h21a == cnt[10:0] ? $signed(32'shada8) : $signed(_GEN_538); // @[FFT.scala 34:12]
  wire [31:0] _GEN_540 = 11'h21b == cnt[10:0] ? $signed(32'shad5e) : $signed(_GEN_539); // @[FFT.scala 34:12]
  wire [31:0] _GEN_541 = 11'h21c == cnt[10:0] ? $signed(32'shad14) : $signed(_GEN_540); // @[FFT.scala 34:12]
  wire [31:0] _GEN_542 = 11'h21d == cnt[10:0] ? $signed(32'shacca) : $signed(_GEN_541); // @[FFT.scala 34:12]
  wire [31:0] _GEN_543 = 11'h21e == cnt[10:0] ? $signed(32'shac80) : $signed(_GEN_542); // @[FFT.scala 34:12]
  wire [31:0] _GEN_544 = 11'h21f == cnt[10:0] ? $signed(32'shac36) : $signed(_GEN_543); // @[FFT.scala 34:12]
  wire [31:0] _GEN_545 = 11'h220 == cnt[10:0] ? $signed(32'shabeb) : $signed(_GEN_544); // @[FFT.scala 34:12]
  wire [31:0] _GEN_546 = 11'h221 == cnt[10:0] ? $signed(32'shaba1) : $signed(_GEN_545); // @[FFT.scala 34:12]
  wire [31:0] _GEN_547 = 11'h222 == cnt[10:0] ? $signed(32'shab56) : $signed(_GEN_546); // @[FFT.scala 34:12]
  wire [31:0] _GEN_548 = 11'h223 == cnt[10:0] ? $signed(32'shab0b) : $signed(_GEN_547); // @[FFT.scala 34:12]
  wire [31:0] _GEN_549 = 11'h224 == cnt[10:0] ? $signed(32'shaac1) : $signed(_GEN_548); // @[FFT.scala 34:12]
  wire [31:0] _GEN_550 = 11'h225 == cnt[10:0] ? $signed(32'shaa76) : $signed(_GEN_549); // @[FFT.scala 34:12]
  wire [31:0] _GEN_551 = 11'h226 == cnt[10:0] ? $signed(32'shaa2a) : $signed(_GEN_550); // @[FFT.scala 34:12]
  wire [31:0] _GEN_552 = 11'h227 == cnt[10:0] ? $signed(32'sha9df) : $signed(_GEN_551); // @[FFT.scala 34:12]
  wire [31:0] _GEN_553 = 11'h228 == cnt[10:0] ? $signed(32'sha994) : $signed(_GEN_552); // @[FFT.scala 34:12]
  wire [31:0] _GEN_554 = 11'h229 == cnt[10:0] ? $signed(32'sha949) : $signed(_GEN_553); // @[FFT.scala 34:12]
  wire [31:0] _GEN_555 = 11'h22a == cnt[10:0] ? $signed(32'sha8fd) : $signed(_GEN_554); // @[FFT.scala 34:12]
  wire [31:0] _GEN_556 = 11'h22b == cnt[10:0] ? $signed(32'sha8b2) : $signed(_GEN_555); // @[FFT.scala 34:12]
  wire [31:0] _GEN_557 = 11'h22c == cnt[10:0] ? $signed(32'sha866) : $signed(_GEN_556); // @[FFT.scala 34:12]
  wire [31:0] _GEN_558 = 11'h22d == cnt[10:0] ? $signed(32'sha81a) : $signed(_GEN_557); // @[FFT.scala 34:12]
  wire [31:0] _GEN_559 = 11'h22e == cnt[10:0] ? $signed(32'sha7ce) : $signed(_GEN_558); // @[FFT.scala 34:12]
  wire [31:0] _GEN_560 = 11'h22f == cnt[10:0] ? $signed(32'sha782) : $signed(_GEN_559); // @[FFT.scala 34:12]
  wire [31:0] _GEN_561 = 11'h230 == cnt[10:0] ? $signed(32'sha736) : $signed(_GEN_560); // @[FFT.scala 34:12]
  wire [31:0] _GEN_562 = 11'h231 == cnt[10:0] ? $signed(32'sha6ea) : $signed(_GEN_561); // @[FFT.scala 34:12]
  wire [31:0] _GEN_563 = 11'h232 == cnt[10:0] ? $signed(32'sha69e) : $signed(_GEN_562); // @[FFT.scala 34:12]
  wire [31:0] _GEN_564 = 11'h233 == cnt[10:0] ? $signed(32'sha652) : $signed(_GEN_563); // @[FFT.scala 34:12]
  wire [31:0] _GEN_565 = 11'h234 == cnt[10:0] ? $signed(32'sha605) : $signed(_GEN_564); // @[FFT.scala 34:12]
  wire [31:0] _GEN_566 = 11'h235 == cnt[10:0] ? $signed(32'sha5b8) : $signed(_GEN_565); // @[FFT.scala 34:12]
  wire [31:0] _GEN_567 = 11'h236 == cnt[10:0] ? $signed(32'sha56c) : $signed(_GEN_566); // @[FFT.scala 34:12]
  wire [31:0] _GEN_568 = 11'h237 == cnt[10:0] ? $signed(32'sha51f) : $signed(_GEN_567); // @[FFT.scala 34:12]
  wire [31:0] _GEN_569 = 11'h238 == cnt[10:0] ? $signed(32'sha4d2) : $signed(_GEN_568); // @[FFT.scala 34:12]
  wire [31:0] _GEN_570 = 11'h239 == cnt[10:0] ? $signed(32'sha485) : $signed(_GEN_569); // @[FFT.scala 34:12]
  wire [31:0] _GEN_571 = 11'h23a == cnt[10:0] ? $signed(32'sha438) : $signed(_GEN_570); // @[FFT.scala 34:12]
  wire [31:0] _GEN_572 = 11'h23b == cnt[10:0] ? $signed(32'sha3eb) : $signed(_GEN_571); // @[FFT.scala 34:12]
  wire [31:0] _GEN_573 = 11'h23c == cnt[10:0] ? $signed(32'sha39e) : $signed(_GEN_572); // @[FFT.scala 34:12]
  wire [31:0] _GEN_574 = 11'h23d == cnt[10:0] ? $signed(32'sha350) : $signed(_GEN_573); // @[FFT.scala 34:12]
  wire [31:0] _GEN_575 = 11'h23e == cnt[10:0] ? $signed(32'sha303) : $signed(_GEN_574); // @[FFT.scala 34:12]
  wire [31:0] _GEN_576 = 11'h23f == cnt[10:0] ? $signed(32'sha2b5) : $signed(_GEN_575); // @[FFT.scala 34:12]
  wire [31:0] _GEN_577 = 11'h240 == cnt[10:0] ? $signed(32'sha268) : $signed(_GEN_576); // @[FFT.scala 34:12]
  wire [31:0] _GEN_578 = 11'h241 == cnt[10:0] ? $signed(32'sha21a) : $signed(_GEN_577); // @[FFT.scala 34:12]
  wire [31:0] _GEN_579 = 11'h242 == cnt[10:0] ? $signed(32'sha1cc) : $signed(_GEN_578); // @[FFT.scala 34:12]
  wire [31:0] _GEN_580 = 11'h243 == cnt[10:0] ? $signed(32'sha17e) : $signed(_GEN_579); // @[FFT.scala 34:12]
  wire [31:0] _GEN_581 = 11'h244 == cnt[10:0] ? $signed(32'sha130) : $signed(_GEN_580); // @[FFT.scala 34:12]
  wire [31:0] _GEN_582 = 11'h245 == cnt[10:0] ? $signed(32'sha0e2) : $signed(_GEN_581); // @[FFT.scala 34:12]
  wire [31:0] _GEN_583 = 11'h246 == cnt[10:0] ? $signed(32'sha094) : $signed(_GEN_582); // @[FFT.scala 34:12]
  wire [31:0] _GEN_584 = 11'h247 == cnt[10:0] ? $signed(32'sha045) : $signed(_GEN_583); // @[FFT.scala 34:12]
  wire [31:0] _GEN_585 = 11'h248 == cnt[10:0] ? $signed(32'sh9ff7) : $signed(_GEN_584); // @[FFT.scala 34:12]
  wire [31:0] _GEN_586 = 11'h249 == cnt[10:0] ? $signed(32'sh9fa8) : $signed(_GEN_585); // @[FFT.scala 34:12]
  wire [31:0] _GEN_587 = 11'h24a == cnt[10:0] ? $signed(32'sh9f5a) : $signed(_GEN_586); // @[FFT.scala 34:12]
  wire [31:0] _GEN_588 = 11'h24b == cnt[10:0] ? $signed(32'sh9f0b) : $signed(_GEN_587); // @[FFT.scala 34:12]
  wire [31:0] _GEN_589 = 11'h24c == cnt[10:0] ? $signed(32'sh9ebc) : $signed(_GEN_588); // @[FFT.scala 34:12]
  wire [31:0] _GEN_590 = 11'h24d == cnt[10:0] ? $signed(32'sh9e6d) : $signed(_GEN_589); // @[FFT.scala 34:12]
  wire [31:0] _GEN_591 = 11'h24e == cnt[10:0] ? $signed(32'sh9e1e) : $signed(_GEN_590); // @[FFT.scala 34:12]
  wire [31:0] _GEN_592 = 11'h24f == cnt[10:0] ? $signed(32'sh9dcf) : $signed(_GEN_591); // @[FFT.scala 34:12]
  wire [31:0] _GEN_593 = 11'h250 == cnt[10:0] ? $signed(32'sh9d80) : $signed(_GEN_592); // @[FFT.scala 34:12]
  wire [31:0] _GEN_594 = 11'h251 == cnt[10:0] ? $signed(32'sh9d31) : $signed(_GEN_593); // @[FFT.scala 34:12]
  wire [31:0] _GEN_595 = 11'h252 == cnt[10:0] ? $signed(32'sh9ce1) : $signed(_GEN_594); // @[FFT.scala 34:12]
  wire [31:0] _GEN_596 = 11'h253 == cnt[10:0] ? $signed(32'sh9c92) : $signed(_GEN_595); // @[FFT.scala 34:12]
  wire [31:0] _GEN_597 = 11'h254 == cnt[10:0] ? $signed(32'sh9c42) : $signed(_GEN_596); // @[FFT.scala 34:12]
  wire [31:0] _GEN_598 = 11'h255 == cnt[10:0] ? $signed(32'sh9bf2) : $signed(_GEN_597); // @[FFT.scala 34:12]
  wire [31:0] _GEN_599 = 11'h256 == cnt[10:0] ? $signed(32'sh9ba3) : $signed(_GEN_598); // @[FFT.scala 34:12]
  wire [31:0] _GEN_600 = 11'h257 == cnt[10:0] ? $signed(32'sh9b53) : $signed(_GEN_599); // @[FFT.scala 34:12]
  wire [31:0] _GEN_601 = 11'h258 == cnt[10:0] ? $signed(32'sh9b03) : $signed(_GEN_600); // @[FFT.scala 34:12]
  wire [31:0] _GEN_602 = 11'h259 == cnt[10:0] ? $signed(32'sh9ab3) : $signed(_GEN_601); // @[FFT.scala 34:12]
  wire [31:0] _GEN_603 = 11'h25a == cnt[10:0] ? $signed(32'sh9a63) : $signed(_GEN_602); // @[FFT.scala 34:12]
  wire [31:0] _GEN_604 = 11'h25b == cnt[10:0] ? $signed(32'sh9a12) : $signed(_GEN_603); // @[FFT.scala 34:12]
  wire [31:0] _GEN_605 = 11'h25c == cnt[10:0] ? $signed(32'sh99c2) : $signed(_GEN_604); // @[FFT.scala 34:12]
  wire [31:0] _GEN_606 = 11'h25d == cnt[10:0] ? $signed(32'sh9972) : $signed(_GEN_605); // @[FFT.scala 34:12]
  wire [31:0] _GEN_607 = 11'h25e == cnt[10:0] ? $signed(32'sh9921) : $signed(_GEN_606); // @[FFT.scala 34:12]
  wire [31:0] _GEN_608 = 11'h25f == cnt[10:0] ? $signed(32'sh98d0) : $signed(_GEN_607); // @[FFT.scala 34:12]
  wire [31:0] _GEN_609 = 11'h260 == cnt[10:0] ? $signed(32'sh9880) : $signed(_GEN_608); // @[FFT.scala 34:12]
  wire [31:0] _GEN_610 = 11'h261 == cnt[10:0] ? $signed(32'sh982f) : $signed(_GEN_609); // @[FFT.scala 34:12]
  wire [31:0] _GEN_611 = 11'h262 == cnt[10:0] ? $signed(32'sh97de) : $signed(_GEN_610); // @[FFT.scala 34:12]
  wire [31:0] _GEN_612 = 11'h263 == cnt[10:0] ? $signed(32'sh978d) : $signed(_GEN_611); // @[FFT.scala 34:12]
  wire [31:0] _GEN_613 = 11'h264 == cnt[10:0] ? $signed(32'sh973c) : $signed(_GEN_612); // @[FFT.scala 34:12]
  wire [31:0] _GEN_614 = 11'h265 == cnt[10:0] ? $signed(32'sh96eb) : $signed(_GEN_613); // @[FFT.scala 34:12]
  wire [31:0] _GEN_615 = 11'h266 == cnt[10:0] ? $signed(32'sh969a) : $signed(_GEN_614); // @[FFT.scala 34:12]
  wire [31:0] _GEN_616 = 11'h267 == cnt[10:0] ? $signed(32'sh9648) : $signed(_GEN_615); // @[FFT.scala 34:12]
  wire [31:0] _GEN_617 = 11'h268 == cnt[10:0] ? $signed(32'sh95f7) : $signed(_GEN_616); // @[FFT.scala 34:12]
  wire [31:0] _GEN_618 = 11'h269 == cnt[10:0] ? $signed(32'sh95a5) : $signed(_GEN_617); // @[FFT.scala 34:12]
  wire [31:0] _GEN_619 = 11'h26a == cnt[10:0] ? $signed(32'sh9554) : $signed(_GEN_618); // @[FFT.scala 34:12]
  wire [31:0] _GEN_620 = 11'h26b == cnt[10:0] ? $signed(32'sh9502) : $signed(_GEN_619); // @[FFT.scala 34:12]
  wire [31:0] _GEN_621 = 11'h26c == cnt[10:0] ? $signed(32'sh94b0) : $signed(_GEN_620); // @[FFT.scala 34:12]
  wire [31:0] _GEN_622 = 11'h26d == cnt[10:0] ? $signed(32'sh945e) : $signed(_GEN_621); // @[FFT.scala 34:12]
  wire [31:0] _GEN_623 = 11'h26e == cnt[10:0] ? $signed(32'sh940c) : $signed(_GEN_622); // @[FFT.scala 34:12]
  wire [31:0] _GEN_624 = 11'h26f == cnt[10:0] ? $signed(32'sh93ba) : $signed(_GEN_623); // @[FFT.scala 34:12]
  wire [31:0] _GEN_625 = 11'h270 == cnt[10:0] ? $signed(32'sh9368) : $signed(_GEN_624); // @[FFT.scala 34:12]
  wire [31:0] _GEN_626 = 11'h271 == cnt[10:0] ? $signed(32'sh9316) : $signed(_GEN_625); // @[FFT.scala 34:12]
  wire [31:0] _GEN_627 = 11'h272 == cnt[10:0] ? $signed(32'sh92c4) : $signed(_GEN_626); // @[FFT.scala 34:12]
  wire [31:0] _GEN_628 = 11'h273 == cnt[10:0] ? $signed(32'sh9271) : $signed(_GEN_627); // @[FFT.scala 34:12]
  wire [31:0] _GEN_629 = 11'h274 == cnt[10:0] ? $signed(32'sh921f) : $signed(_GEN_628); // @[FFT.scala 34:12]
  wire [31:0] _GEN_630 = 11'h275 == cnt[10:0] ? $signed(32'sh91cc) : $signed(_GEN_629); // @[FFT.scala 34:12]
  wire [31:0] _GEN_631 = 11'h276 == cnt[10:0] ? $signed(32'sh9179) : $signed(_GEN_630); // @[FFT.scala 34:12]
  wire [31:0] _GEN_632 = 11'h277 == cnt[10:0] ? $signed(32'sh9127) : $signed(_GEN_631); // @[FFT.scala 34:12]
  wire [31:0] _GEN_633 = 11'h278 == cnt[10:0] ? $signed(32'sh90d4) : $signed(_GEN_632); // @[FFT.scala 34:12]
  wire [31:0] _GEN_634 = 11'h279 == cnt[10:0] ? $signed(32'sh9081) : $signed(_GEN_633); // @[FFT.scala 34:12]
  wire [31:0] _GEN_635 = 11'h27a == cnt[10:0] ? $signed(32'sh902e) : $signed(_GEN_634); // @[FFT.scala 34:12]
  wire [31:0] _GEN_636 = 11'h27b == cnt[10:0] ? $signed(32'sh8fdb) : $signed(_GEN_635); // @[FFT.scala 34:12]
  wire [31:0] _GEN_637 = 11'h27c == cnt[10:0] ? $signed(32'sh8f88) : $signed(_GEN_636); // @[FFT.scala 34:12]
  wire [31:0] _GEN_638 = 11'h27d == cnt[10:0] ? $signed(32'sh8f34) : $signed(_GEN_637); // @[FFT.scala 34:12]
  wire [31:0] _GEN_639 = 11'h27e == cnt[10:0] ? $signed(32'sh8ee1) : $signed(_GEN_638); // @[FFT.scala 34:12]
  wire [31:0] _GEN_640 = 11'h27f == cnt[10:0] ? $signed(32'sh8e8d) : $signed(_GEN_639); // @[FFT.scala 34:12]
  wire [31:0] _GEN_641 = 11'h280 == cnt[10:0] ? $signed(32'sh8e3a) : $signed(_GEN_640); // @[FFT.scala 34:12]
  wire [31:0] _GEN_642 = 11'h281 == cnt[10:0] ? $signed(32'sh8de6) : $signed(_GEN_641); // @[FFT.scala 34:12]
  wire [31:0] _GEN_643 = 11'h282 == cnt[10:0] ? $signed(32'sh8d93) : $signed(_GEN_642); // @[FFT.scala 34:12]
  wire [31:0] _GEN_644 = 11'h283 == cnt[10:0] ? $signed(32'sh8d3f) : $signed(_GEN_643); // @[FFT.scala 34:12]
  wire [31:0] _GEN_645 = 11'h284 == cnt[10:0] ? $signed(32'sh8ceb) : $signed(_GEN_644); // @[FFT.scala 34:12]
  wire [31:0] _GEN_646 = 11'h285 == cnt[10:0] ? $signed(32'sh8c97) : $signed(_GEN_645); // @[FFT.scala 34:12]
  wire [31:0] _GEN_647 = 11'h286 == cnt[10:0] ? $signed(32'sh8c43) : $signed(_GEN_646); // @[FFT.scala 34:12]
  wire [31:0] _GEN_648 = 11'h287 == cnt[10:0] ? $signed(32'sh8bef) : $signed(_GEN_647); // @[FFT.scala 34:12]
  wire [31:0] _GEN_649 = 11'h288 == cnt[10:0] ? $signed(32'sh8b9a) : $signed(_GEN_648); // @[FFT.scala 34:12]
  wire [31:0] _GEN_650 = 11'h289 == cnt[10:0] ? $signed(32'sh8b46) : $signed(_GEN_649); // @[FFT.scala 34:12]
  wire [31:0] _GEN_651 = 11'h28a == cnt[10:0] ? $signed(32'sh8af2) : $signed(_GEN_650); // @[FFT.scala 34:12]
  wire [31:0] _GEN_652 = 11'h28b == cnt[10:0] ? $signed(32'sh8a9d) : $signed(_GEN_651); // @[FFT.scala 34:12]
  wire [31:0] _GEN_653 = 11'h28c == cnt[10:0] ? $signed(32'sh8a49) : $signed(_GEN_652); // @[FFT.scala 34:12]
  wire [31:0] _GEN_654 = 11'h28d == cnt[10:0] ? $signed(32'sh89f4) : $signed(_GEN_653); // @[FFT.scala 34:12]
  wire [31:0] _GEN_655 = 11'h28e == cnt[10:0] ? $signed(32'sh899f) : $signed(_GEN_654); // @[FFT.scala 34:12]
  wire [31:0] _GEN_656 = 11'h28f == cnt[10:0] ? $signed(32'sh894a) : $signed(_GEN_655); // @[FFT.scala 34:12]
  wire [31:0] _GEN_657 = 11'h290 == cnt[10:0] ? $signed(32'sh88f6) : $signed(_GEN_656); // @[FFT.scala 34:12]
  wire [31:0] _GEN_658 = 11'h291 == cnt[10:0] ? $signed(32'sh88a1) : $signed(_GEN_657); // @[FFT.scala 34:12]
  wire [31:0] _GEN_659 = 11'h292 == cnt[10:0] ? $signed(32'sh884c) : $signed(_GEN_658); // @[FFT.scala 34:12]
  wire [31:0] _GEN_660 = 11'h293 == cnt[10:0] ? $signed(32'sh87f6) : $signed(_GEN_659); // @[FFT.scala 34:12]
  wire [31:0] _GEN_661 = 11'h294 == cnt[10:0] ? $signed(32'sh87a1) : $signed(_GEN_660); // @[FFT.scala 34:12]
  wire [31:0] _GEN_662 = 11'h295 == cnt[10:0] ? $signed(32'sh874c) : $signed(_GEN_661); // @[FFT.scala 34:12]
  wire [31:0] _GEN_663 = 11'h296 == cnt[10:0] ? $signed(32'sh86f7) : $signed(_GEN_662); // @[FFT.scala 34:12]
  wire [31:0] _GEN_664 = 11'h297 == cnt[10:0] ? $signed(32'sh86a1) : $signed(_GEN_663); // @[FFT.scala 34:12]
  wire [31:0] _GEN_665 = 11'h298 == cnt[10:0] ? $signed(32'sh864c) : $signed(_GEN_664); // @[FFT.scala 34:12]
  wire [31:0] _GEN_666 = 11'h299 == cnt[10:0] ? $signed(32'sh85f6) : $signed(_GEN_665); // @[FFT.scala 34:12]
  wire [31:0] _GEN_667 = 11'h29a == cnt[10:0] ? $signed(32'sh85a0) : $signed(_GEN_666); // @[FFT.scala 34:12]
  wire [31:0] _GEN_668 = 11'h29b == cnt[10:0] ? $signed(32'sh854a) : $signed(_GEN_667); // @[FFT.scala 34:12]
  wire [31:0] _GEN_669 = 11'h29c == cnt[10:0] ? $signed(32'sh84f5) : $signed(_GEN_668); // @[FFT.scala 34:12]
  wire [31:0] _GEN_670 = 11'h29d == cnt[10:0] ? $signed(32'sh849f) : $signed(_GEN_669); // @[FFT.scala 34:12]
  wire [31:0] _GEN_671 = 11'h29e == cnt[10:0] ? $signed(32'sh8449) : $signed(_GEN_670); // @[FFT.scala 34:12]
  wire [31:0] _GEN_672 = 11'h29f == cnt[10:0] ? $signed(32'sh83f2) : $signed(_GEN_671); // @[FFT.scala 34:12]
  wire [31:0] _GEN_673 = 11'h2a0 == cnt[10:0] ? $signed(32'sh839c) : $signed(_GEN_672); // @[FFT.scala 34:12]
  wire [31:0] _GEN_674 = 11'h2a1 == cnt[10:0] ? $signed(32'sh8346) : $signed(_GEN_673); // @[FFT.scala 34:12]
  wire [31:0] _GEN_675 = 11'h2a2 == cnt[10:0] ? $signed(32'sh82f0) : $signed(_GEN_674); // @[FFT.scala 34:12]
  wire [31:0] _GEN_676 = 11'h2a3 == cnt[10:0] ? $signed(32'sh8299) : $signed(_GEN_675); // @[FFT.scala 34:12]
  wire [31:0] _GEN_677 = 11'h2a4 == cnt[10:0] ? $signed(32'sh8243) : $signed(_GEN_676); // @[FFT.scala 34:12]
  wire [31:0] _GEN_678 = 11'h2a5 == cnt[10:0] ? $signed(32'sh81ec) : $signed(_GEN_677); // @[FFT.scala 34:12]
  wire [31:0] _GEN_679 = 11'h2a6 == cnt[10:0] ? $signed(32'sh8195) : $signed(_GEN_678); // @[FFT.scala 34:12]
  wire [31:0] _GEN_680 = 11'h2a7 == cnt[10:0] ? $signed(32'sh813f) : $signed(_GEN_679); // @[FFT.scala 34:12]
  wire [31:0] _GEN_681 = 11'h2a8 == cnt[10:0] ? $signed(32'sh80e8) : $signed(_GEN_680); // @[FFT.scala 34:12]
  wire [31:0] _GEN_682 = 11'h2a9 == cnt[10:0] ? $signed(32'sh8091) : $signed(_GEN_681); // @[FFT.scala 34:12]
  wire [31:0] _GEN_683 = 11'h2aa == cnt[10:0] ? $signed(32'sh803a) : $signed(_GEN_682); // @[FFT.scala 34:12]
  wire [31:0] _GEN_684 = 11'h2ab == cnt[10:0] ? $signed(32'sh7fe3) : $signed(_GEN_683); // @[FFT.scala 34:12]
  wire [31:0] _GEN_685 = 11'h2ac == cnt[10:0] ? $signed(32'sh7f8c) : $signed(_GEN_684); // @[FFT.scala 34:12]
  wire [31:0] _GEN_686 = 11'h2ad == cnt[10:0] ? $signed(32'sh7f35) : $signed(_GEN_685); // @[FFT.scala 34:12]
  wire [31:0] _GEN_687 = 11'h2ae == cnt[10:0] ? $signed(32'sh7edd) : $signed(_GEN_686); // @[FFT.scala 34:12]
  wire [31:0] _GEN_688 = 11'h2af == cnt[10:0] ? $signed(32'sh7e86) : $signed(_GEN_687); // @[FFT.scala 34:12]
  wire [31:0] _GEN_689 = 11'h2b0 == cnt[10:0] ? $signed(32'sh7e2f) : $signed(_GEN_688); // @[FFT.scala 34:12]
  wire [31:0] _GEN_690 = 11'h2b1 == cnt[10:0] ? $signed(32'sh7dd7) : $signed(_GEN_689); // @[FFT.scala 34:12]
  wire [31:0] _GEN_691 = 11'h2b2 == cnt[10:0] ? $signed(32'sh7d7f) : $signed(_GEN_690); // @[FFT.scala 34:12]
  wire [31:0] _GEN_692 = 11'h2b3 == cnt[10:0] ? $signed(32'sh7d28) : $signed(_GEN_691); // @[FFT.scala 34:12]
  wire [31:0] _GEN_693 = 11'h2b4 == cnt[10:0] ? $signed(32'sh7cd0) : $signed(_GEN_692); // @[FFT.scala 34:12]
  wire [31:0] _GEN_694 = 11'h2b5 == cnt[10:0] ? $signed(32'sh7c78) : $signed(_GEN_693); // @[FFT.scala 34:12]
  wire [31:0] _GEN_695 = 11'h2b6 == cnt[10:0] ? $signed(32'sh7c20) : $signed(_GEN_694); // @[FFT.scala 34:12]
  wire [31:0] _GEN_696 = 11'h2b7 == cnt[10:0] ? $signed(32'sh7bc8) : $signed(_GEN_695); // @[FFT.scala 34:12]
  wire [31:0] _GEN_697 = 11'h2b8 == cnt[10:0] ? $signed(32'sh7b70) : $signed(_GEN_696); // @[FFT.scala 34:12]
  wire [31:0] _GEN_698 = 11'h2b9 == cnt[10:0] ? $signed(32'sh7b18) : $signed(_GEN_697); // @[FFT.scala 34:12]
  wire [31:0] _GEN_699 = 11'h2ba == cnt[10:0] ? $signed(32'sh7ac0) : $signed(_GEN_698); // @[FFT.scala 34:12]
  wire [31:0] _GEN_700 = 11'h2bb == cnt[10:0] ? $signed(32'sh7a68) : $signed(_GEN_699); // @[FFT.scala 34:12]
  wire [31:0] _GEN_701 = 11'h2bc == cnt[10:0] ? $signed(32'sh7a10) : $signed(_GEN_700); // @[FFT.scala 34:12]
  wire [31:0] _GEN_702 = 11'h2bd == cnt[10:0] ? $signed(32'sh79b7) : $signed(_GEN_701); // @[FFT.scala 34:12]
  wire [31:0] _GEN_703 = 11'h2be == cnt[10:0] ? $signed(32'sh795f) : $signed(_GEN_702); // @[FFT.scala 34:12]
  wire [31:0] _GEN_704 = 11'h2bf == cnt[10:0] ? $signed(32'sh7906) : $signed(_GEN_703); // @[FFT.scala 34:12]
  wire [31:0] _GEN_705 = 11'h2c0 == cnt[10:0] ? $signed(32'sh78ad) : $signed(_GEN_704); // @[FFT.scala 34:12]
  wire [31:0] _GEN_706 = 11'h2c1 == cnt[10:0] ? $signed(32'sh7855) : $signed(_GEN_705); // @[FFT.scala 34:12]
  wire [31:0] _GEN_707 = 11'h2c2 == cnt[10:0] ? $signed(32'sh77fc) : $signed(_GEN_706); // @[FFT.scala 34:12]
  wire [31:0] _GEN_708 = 11'h2c3 == cnt[10:0] ? $signed(32'sh77a3) : $signed(_GEN_707); // @[FFT.scala 34:12]
  wire [31:0] _GEN_709 = 11'h2c4 == cnt[10:0] ? $signed(32'sh774a) : $signed(_GEN_708); // @[FFT.scala 34:12]
  wire [31:0] _GEN_710 = 11'h2c5 == cnt[10:0] ? $signed(32'sh76f1) : $signed(_GEN_709); // @[FFT.scala 34:12]
  wire [31:0] _GEN_711 = 11'h2c6 == cnt[10:0] ? $signed(32'sh7698) : $signed(_GEN_710); // @[FFT.scala 34:12]
  wire [31:0] _GEN_712 = 11'h2c7 == cnt[10:0] ? $signed(32'sh763f) : $signed(_GEN_711); // @[FFT.scala 34:12]
  wire [31:0] _GEN_713 = 11'h2c8 == cnt[10:0] ? $signed(32'sh75e6) : $signed(_GEN_712); // @[FFT.scala 34:12]
  wire [31:0] _GEN_714 = 11'h2c9 == cnt[10:0] ? $signed(32'sh758d) : $signed(_GEN_713); // @[FFT.scala 34:12]
  wire [31:0] _GEN_715 = 11'h2ca == cnt[10:0] ? $signed(32'sh7533) : $signed(_GEN_714); // @[FFT.scala 34:12]
  wire [31:0] _GEN_716 = 11'h2cb == cnt[10:0] ? $signed(32'sh74da) : $signed(_GEN_715); // @[FFT.scala 34:12]
  wire [31:0] _GEN_717 = 11'h2cc == cnt[10:0] ? $signed(32'sh7480) : $signed(_GEN_716); // @[FFT.scala 34:12]
  wire [31:0] _GEN_718 = 11'h2cd == cnt[10:0] ? $signed(32'sh7427) : $signed(_GEN_717); // @[FFT.scala 34:12]
  wire [31:0] _GEN_719 = 11'h2ce == cnt[10:0] ? $signed(32'sh73cd) : $signed(_GEN_718); // @[FFT.scala 34:12]
  wire [31:0] _GEN_720 = 11'h2cf == cnt[10:0] ? $signed(32'sh7373) : $signed(_GEN_719); // @[FFT.scala 34:12]
  wire [31:0] _GEN_721 = 11'h2d0 == cnt[10:0] ? $signed(32'sh731a) : $signed(_GEN_720); // @[FFT.scala 34:12]
  wire [31:0] _GEN_722 = 11'h2d1 == cnt[10:0] ? $signed(32'sh72c0) : $signed(_GEN_721); // @[FFT.scala 34:12]
  wire [31:0] _GEN_723 = 11'h2d2 == cnt[10:0] ? $signed(32'sh7266) : $signed(_GEN_722); // @[FFT.scala 34:12]
  wire [31:0] _GEN_724 = 11'h2d3 == cnt[10:0] ? $signed(32'sh720c) : $signed(_GEN_723); // @[FFT.scala 34:12]
  wire [31:0] _GEN_725 = 11'h2d4 == cnt[10:0] ? $signed(32'sh71b2) : $signed(_GEN_724); // @[FFT.scala 34:12]
  wire [31:0] _GEN_726 = 11'h2d5 == cnt[10:0] ? $signed(32'sh7158) : $signed(_GEN_725); // @[FFT.scala 34:12]
  wire [31:0] _GEN_727 = 11'h2d6 == cnt[10:0] ? $signed(32'sh70fe) : $signed(_GEN_726); // @[FFT.scala 34:12]
  wire [31:0] _GEN_728 = 11'h2d7 == cnt[10:0] ? $signed(32'sh70a3) : $signed(_GEN_727); // @[FFT.scala 34:12]
  wire [31:0] _GEN_729 = 11'h2d8 == cnt[10:0] ? $signed(32'sh7049) : $signed(_GEN_728); // @[FFT.scala 34:12]
  wire [31:0] _GEN_730 = 11'h2d9 == cnt[10:0] ? $signed(32'sh6fef) : $signed(_GEN_729); // @[FFT.scala 34:12]
  wire [31:0] _GEN_731 = 11'h2da == cnt[10:0] ? $signed(32'sh6f94) : $signed(_GEN_730); // @[FFT.scala 34:12]
  wire [31:0] _GEN_732 = 11'h2db == cnt[10:0] ? $signed(32'sh6f3a) : $signed(_GEN_731); // @[FFT.scala 34:12]
  wire [31:0] _GEN_733 = 11'h2dc == cnt[10:0] ? $signed(32'sh6edf) : $signed(_GEN_732); // @[FFT.scala 34:12]
  wire [31:0] _GEN_734 = 11'h2dd == cnt[10:0] ? $signed(32'sh6e85) : $signed(_GEN_733); // @[FFT.scala 34:12]
  wire [31:0] _GEN_735 = 11'h2de == cnt[10:0] ? $signed(32'sh6e2a) : $signed(_GEN_734); // @[FFT.scala 34:12]
  wire [31:0] _GEN_736 = 11'h2df == cnt[10:0] ? $signed(32'sh6dcf) : $signed(_GEN_735); // @[FFT.scala 34:12]
  wire [31:0] _GEN_737 = 11'h2e0 == cnt[10:0] ? $signed(32'sh6d74) : $signed(_GEN_736); // @[FFT.scala 34:12]
  wire [31:0] _GEN_738 = 11'h2e1 == cnt[10:0] ? $signed(32'sh6d19) : $signed(_GEN_737); // @[FFT.scala 34:12]
  wire [31:0] _GEN_739 = 11'h2e2 == cnt[10:0] ? $signed(32'sh6cbe) : $signed(_GEN_738); // @[FFT.scala 34:12]
  wire [31:0] _GEN_740 = 11'h2e3 == cnt[10:0] ? $signed(32'sh6c63) : $signed(_GEN_739); // @[FFT.scala 34:12]
  wire [31:0] _GEN_741 = 11'h2e4 == cnt[10:0] ? $signed(32'sh6c08) : $signed(_GEN_740); // @[FFT.scala 34:12]
  wire [31:0] _GEN_742 = 11'h2e5 == cnt[10:0] ? $signed(32'sh6bad) : $signed(_GEN_741); // @[FFT.scala 34:12]
  wire [31:0] _GEN_743 = 11'h2e6 == cnt[10:0] ? $signed(32'sh6b52) : $signed(_GEN_742); // @[FFT.scala 34:12]
  wire [31:0] _GEN_744 = 11'h2e7 == cnt[10:0] ? $signed(32'sh6af6) : $signed(_GEN_743); // @[FFT.scala 34:12]
  wire [31:0] _GEN_745 = 11'h2e8 == cnt[10:0] ? $signed(32'sh6a9b) : $signed(_GEN_744); // @[FFT.scala 34:12]
  wire [31:0] _GEN_746 = 11'h2e9 == cnt[10:0] ? $signed(32'sh6a40) : $signed(_GEN_745); // @[FFT.scala 34:12]
  wire [31:0] _GEN_747 = 11'h2ea == cnt[10:0] ? $signed(32'sh69e4) : $signed(_GEN_746); // @[FFT.scala 34:12]
  wire [31:0] _GEN_748 = 11'h2eb == cnt[10:0] ? $signed(32'sh6989) : $signed(_GEN_747); // @[FFT.scala 34:12]
  wire [31:0] _GEN_749 = 11'h2ec == cnt[10:0] ? $signed(32'sh692d) : $signed(_GEN_748); // @[FFT.scala 34:12]
  wire [31:0] _GEN_750 = 11'h2ed == cnt[10:0] ? $signed(32'sh68d1) : $signed(_GEN_749); // @[FFT.scala 34:12]
  wire [31:0] _GEN_751 = 11'h2ee == cnt[10:0] ? $signed(32'sh6876) : $signed(_GEN_750); // @[FFT.scala 34:12]
  wire [31:0] _GEN_752 = 11'h2ef == cnt[10:0] ? $signed(32'sh681a) : $signed(_GEN_751); // @[FFT.scala 34:12]
  wire [31:0] _GEN_753 = 11'h2f0 == cnt[10:0] ? $signed(32'sh67be) : $signed(_GEN_752); // @[FFT.scala 34:12]
  wire [31:0] _GEN_754 = 11'h2f1 == cnt[10:0] ? $signed(32'sh6762) : $signed(_GEN_753); // @[FFT.scala 34:12]
  wire [31:0] _GEN_755 = 11'h2f2 == cnt[10:0] ? $signed(32'sh6706) : $signed(_GEN_754); // @[FFT.scala 34:12]
  wire [31:0] _GEN_756 = 11'h2f3 == cnt[10:0] ? $signed(32'sh66aa) : $signed(_GEN_755); // @[FFT.scala 34:12]
  wire [31:0] _GEN_757 = 11'h2f4 == cnt[10:0] ? $signed(32'sh664e) : $signed(_GEN_756); // @[FFT.scala 34:12]
  wire [31:0] _GEN_758 = 11'h2f5 == cnt[10:0] ? $signed(32'sh65f2) : $signed(_GEN_757); // @[FFT.scala 34:12]
  wire [31:0] _GEN_759 = 11'h2f6 == cnt[10:0] ? $signed(32'sh6595) : $signed(_GEN_758); // @[FFT.scala 34:12]
  wire [31:0] _GEN_760 = 11'h2f7 == cnt[10:0] ? $signed(32'sh6539) : $signed(_GEN_759); // @[FFT.scala 34:12]
  wire [31:0] _GEN_761 = 11'h2f8 == cnt[10:0] ? $signed(32'sh64dd) : $signed(_GEN_760); // @[FFT.scala 34:12]
  wire [31:0] _GEN_762 = 11'h2f9 == cnt[10:0] ? $signed(32'sh6480) : $signed(_GEN_761); // @[FFT.scala 34:12]
  wire [31:0] _GEN_763 = 11'h2fa == cnt[10:0] ? $signed(32'sh6424) : $signed(_GEN_762); // @[FFT.scala 34:12]
  wire [31:0] _GEN_764 = 11'h2fb == cnt[10:0] ? $signed(32'sh63c7) : $signed(_GEN_763); // @[FFT.scala 34:12]
  wire [31:0] _GEN_765 = 11'h2fc == cnt[10:0] ? $signed(32'sh636b) : $signed(_GEN_764); // @[FFT.scala 34:12]
  wire [31:0] _GEN_766 = 11'h2fd == cnt[10:0] ? $signed(32'sh630e) : $signed(_GEN_765); // @[FFT.scala 34:12]
  wire [31:0] _GEN_767 = 11'h2fe == cnt[10:0] ? $signed(32'sh62b1) : $signed(_GEN_766); // @[FFT.scala 34:12]
  wire [31:0] _GEN_768 = 11'h2ff == cnt[10:0] ? $signed(32'sh6254) : $signed(_GEN_767); // @[FFT.scala 34:12]
  wire [31:0] _GEN_769 = 11'h300 == cnt[10:0] ? $signed(32'sh61f8) : $signed(_GEN_768); // @[FFT.scala 34:12]
  wire [31:0] _GEN_770 = 11'h301 == cnt[10:0] ? $signed(32'sh619b) : $signed(_GEN_769); // @[FFT.scala 34:12]
  wire [31:0] _GEN_771 = 11'h302 == cnt[10:0] ? $signed(32'sh613e) : $signed(_GEN_770); // @[FFT.scala 34:12]
  wire [31:0] _GEN_772 = 11'h303 == cnt[10:0] ? $signed(32'sh60e1) : $signed(_GEN_771); // @[FFT.scala 34:12]
  wire [31:0] _GEN_773 = 11'h304 == cnt[10:0] ? $signed(32'sh6084) : $signed(_GEN_772); // @[FFT.scala 34:12]
  wire [31:0] _GEN_774 = 11'h305 == cnt[10:0] ? $signed(32'sh6026) : $signed(_GEN_773); // @[FFT.scala 34:12]
  wire [31:0] _GEN_775 = 11'h306 == cnt[10:0] ? $signed(32'sh5fc9) : $signed(_GEN_774); // @[FFT.scala 34:12]
  wire [31:0] _GEN_776 = 11'h307 == cnt[10:0] ? $signed(32'sh5f6c) : $signed(_GEN_775); // @[FFT.scala 34:12]
  wire [31:0] _GEN_777 = 11'h308 == cnt[10:0] ? $signed(32'sh5f0f) : $signed(_GEN_776); // @[FFT.scala 34:12]
  wire [31:0] _GEN_778 = 11'h309 == cnt[10:0] ? $signed(32'sh5eb1) : $signed(_GEN_777); // @[FFT.scala 34:12]
  wire [31:0] _GEN_779 = 11'h30a == cnt[10:0] ? $signed(32'sh5e54) : $signed(_GEN_778); // @[FFT.scala 34:12]
  wire [31:0] _GEN_780 = 11'h30b == cnt[10:0] ? $signed(32'sh5df6) : $signed(_GEN_779); // @[FFT.scala 34:12]
  wire [31:0] _GEN_781 = 11'h30c == cnt[10:0] ? $signed(32'sh5d99) : $signed(_GEN_780); // @[FFT.scala 34:12]
  wire [31:0] _GEN_782 = 11'h30d == cnt[10:0] ? $signed(32'sh5d3b) : $signed(_GEN_781); // @[FFT.scala 34:12]
  wire [31:0] _GEN_783 = 11'h30e == cnt[10:0] ? $signed(32'sh5cde) : $signed(_GEN_782); // @[FFT.scala 34:12]
  wire [31:0] _GEN_784 = 11'h30f == cnt[10:0] ? $signed(32'sh5c80) : $signed(_GEN_783); // @[FFT.scala 34:12]
  wire [31:0] _GEN_785 = 11'h310 == cnt[10:0] ? $signed(32'sh5c22) : $signed(_GEN_784); // @[FFT.scala 34:12]
  wire [31:0] _GEN_786 = 11'h311 == cnt[10:0] ? $signed(32'sh5bc4) : $signed(_GEN_785); // @[FFT.scala 34:12]
  wire [31:0] _GEN_787 = 11'h312 == cnt[10:0] ? $signed(32'sh5b66) : $signed(_GEN_786); // @[FFT.scala 34:12]
  wire [31:0] _GEN_788 = 11'h313 == cnt[10:0] ? $signed(32'sh5b08) : $signed(_GEN_787); // @[FFT.scala 34:12]
  wire [31:0] _GEN_789 = 11'h314 == cnt[10:0] ? $signed(32'sh5aaa) : $signed(_GEN_788); // @[FFT.scala 34:12]
  wire [31:0] _GEN_790 = 11'h315 == cnt[10:0] ? $signed(32'sh5a4c) : $signed(_GEN_789); // @[FFT.scala 34:12]
  wire [31:0] _GEN_791 = 11'h316 == cnt[10:0] ? $signed(32'sh59ee) : $signed(_GEN_790); // @[FFT.scala 34:12]
  wire [31:0] _GEN_792 = 11'h317 == cnt[10:0] ? $signed(32'sh5990) : $signed(_GEN_791); // @[FFT.scala 34:12]
  wire [31:0] _GEN_793 = 11'h318 == cnt[10:0] ? $signed(32'sh5932) : $signed(_GEN_792); // @[FFT.scala 34:12]
  wire [31:0] _GEN_794 = 11'h319 == cnt[10:0] ? $signed(32'sh58d4) : $signed(_GEN_793); // @[FFT.scala 34:12]
  wire [31:0] _GEN_795 = 11'h31a == cnt[10:0] ? $signed(32'sh5875) : $signed(_GEN_794); // @[FFT.scala 34:12]
  wire [31:0] _GEN_796 = 11'h31b == cnt[10:0] ? $signed(32'sh5817) : $signed(_GEN_795); // @[FFT.scala 34:12]
  wire [31:0] _GEN_797 = 11'h31c == cnt[10:0] ? $signed(32'sh57b9) : $signed(_GEN_796); // @[FFT.scala 34:12]
  wire [31:0] _GEN_798 = 11'h31d == cnt[10:0] ? $signed(32'sh575a) : $signed(_GEN_797); // @[FFT.scala 34:12]
  wire [31:0] _GEN_799 = 11'h31e == cnt[10:0] ? $signed(32'sh56fc) : $signed(_GEN_798); // @[FFT.scala 34:12]
  wire [31:0] _GEN_800 = 11'h31f == cnt[10:0] ? $signed(32'sh569d) : $signed(_GEN_799); // @[FFT.scala 34:12]
  wire [31:0] _GEN_801 = 11'h320 == cnt[10:0] ? $signed(32'sh563e) : $signed(_GEN_800); // @[FFT.scala 34:12]
  wire [31:0] _GEN_802 = 11'h321 == cnt[10:0] ? $signed(32'sh55e0) : $signed(_GEN_801); // @[FFT.scala 34:12]
  wire [31:0] _GEN_803 = 11'h322 == cnt[10:0] ? $signed(32'sh5581) : $signed(_GEN_802); // @[FFT.scala 34:12]
  wire [31:0] _GEN_804 = 11'h323 == cnt[10:0] ? $signed(32'sh5522) : $signed(_GEN_803); // @[FFT.scala 34:12]
  wire [31:0] _GEN_805 = 11'h324 == cnt[10:0] ? $signed(32'sh54c3) : $signed(_GEN_804); // @[FFT.scala 34:12]
  wire [31:0] _GEN_806 = 11'h325 == cnt[10:0] ? $signed(32'sh5464) : $signed(_GEN_805); // @[FFT.scala 34:12]
  wire [31:0] _GEN_807 = 11'h326 == cnt[10:0] ? $signed(32'sh5406) : $signed(_GEN_806); // @[FFT.scala 34:12]
  wire [31:0] _GEN_808 = 11'h327 == cnt[10:0] ? $signed(32'sh53a7) : $signed(_GEN_807); // @[FFT.scala 34:12]
  wire [31:0] _GEN_809 = 11'h328 == cnt[10:0] ? $signed(32'sh5348) : $signed(_GEN_808); // @[FFT.scala 34:12]
  wire [31:0] _GEN_810 = 11'h329 == cnt[10:0] ? $signed(32'sh52e8) : $signed(_GEN_809); // @[FFT.scala 34:12]
  wire [31:0] _GEN_811 = 11'h32a == cnt[10:0] ? $signed(32'sh5289) : $signed(_GEN_810); // @[FFT.scala 34:12]
  wire [31:0] _GEN_812 = 11'h32b == cnt[10:0] ? $signed(32'sh522a) : $signed(_GEN_811); // @[FFT.scala 34:12]
  wire [31:0] _GEN_813 = 11'h32c == cnt[10:0] ? $signed(32'sh51cb) : $signed(_GEN_812); // @[FFT.scala 34:12]
  wire [31:0] _GEN_814 = 11'h32d == cnt[10:0] ? $signed(32'sh516c) : $signed(_GEN_813); // @[FFT.scala 34:12]
  wire [31:0] _GEN_815 = 11'h32e == cnt[10:0] ? $signed(32'sh510c) : $signed(_GEN_814); // @[FFT.scala 34:12]
  wire [31:0] _GEN_816 = 11'h32f == cnt[10:0] ? $signed(32'sh50ad) : $signed(_GEN_815); // @[FFT.scala 34:12]
  wire [31:0] _GEN_817 = 11'h330 == cnt[10:0] ? $signed(32'sh504d) : $signed(_GEN_816); // @[FFT.scala 34:12]
  wire [31:0] _GEN_818 = 11'h331 == cnt[10:0] ? $signed(32'sh4fee) : $signed(_GEN_817); // @[FFT.scala 34:12]
  wire [31:0] _GEN_819 = 11'h332 == cnt[10:0] ? $signed(32'sh4f8e) : $signed(_GEN_818); // @[FFT.scala 34:12]
  wire [31:0] _GEN_820 = 11'h333 == cnt[10:0] ? $signed(32'sh4f2f) : $signed(_GEN_819); // @[FFT.scala 34:12]
  wire [31:0] _GEN_821 = 11'h334 == cnt[10:0] ? $signed(32'sh4ecf) : $signed(_GEN_820); // @[FFT.scala 34:12]
  wire [31:0] _GEN_822 = 11'h335 == cnt[10:0] ? $signed(32'sh4e70) : $signed(_GEN_821); // @[FFT.scala 34:12]
  wire [31:0] _GEN_823 = 11'h336 == cnt[10:0] ? $signed(32'sh4e10) : $signed(_GEN_822); // @[FFT.scala 34:12]
  wire [31:0] _GEN_824 = 11'h337 == cnt[10:0] ? $signed(32'sh4db0) : $signed(_GEN_823); // @[FFT.scala 34:12]
  wire [31:0] _GEN_825 = 11'h338 == cnt[10:0] ? $signed(32'sh4d50) : $signed(_GEN_824); // @[FFT.scala 34:12]
  wire [31:0] _GEN_826 = 11'h339 == cnt[10:0] ? $signed(32'sh4cf0) : $signed(_GEN_825); // @[FFT.scala 34:12]
  wire [31:0] _GEN_827 = 11'h33a == cnt[10:0] ? $signed(32'sh4c90) : $signed(_GEN_826); // @[FFT.scala 34:12]
  wire [31:0] _GEN_828 = 11'h33b == cnt[10:0] ? $signed(32'sh4c31) : $signed(_GEN_827); // @[FFT.scala 34:12]
  wire [31:0] _GEN_829 = 11'h33c == cnt[10:0] ? $signed(32'sh4bd1) : $signed(_GEN_828); // @[FFT.scala 34:12]
  wire [31:0] _GEN_830 = 11'h33d == cnt[10:0] ? $signed(32'sh4b71) : $signed(_GEN_829); // @[FFT.scala 34:12]
  wire [31:0] _GEN_831 = 11'h33e == cnt[10:0] ? $signed(32'sh4b10) : $signed(_GEN_830); // @[FFT.scala 34:12]
  wire [31:0] _GEN_832 = 11'h33f == cnt[10:0] ? $signed(32'sh4ab0) : $signed(_GEN_831); // @[FFT.scala 34:12]
  wire [31:0] _GEN_833 = 11'h340 == cnt[10:0] ? $signed(32'sh4a50) : $signed(_GEN_832); // @[FFT.scala 34:12]
  wire [31:0] _GEN_834 = 11'h341 == cnt[10:0] ? $signed(32'sh49f0) : $signed(_GEN_833); // @[FFT.scala 34:12]
  wire [31:0] _GEN_835 = 11'h342 == cnt[10:0] ? $signed(32'sh4990) : $signed(_GEN_834); // @[FFT.scala 34:12]
  wire [31:0] _GEN_836 = 11'h343 == cnt[10:0] ? $signed(32'sh492f) : $signed(_GEN_835); // @[FFT.scala 34:12]
  wire [31:0] _GEN_837 = 11'h344 == cnt[10:0] ? $signed(32'sh48cf) : $signed(_GEN_836); // @[FFT.scala 34:12]
  wire [31:0] _GEN_838 = 11'h345 == cnt[10:0] ? $signed(32'sh486f) : $signed(_GEN_837); // @[FFT.scala 34:12]
  wire [31:0] _GEN_839 = 11'h346 == cnt[10:0] ? $signed(32'sh480e) : $signed(_GEN_838); // @[FFT.scala 34:12]
  wire [31:0] _GEN_840 = 11'h347 == cnt[10:0] ? $signed(32'sh47ae) : $signed(_GEN_839); // @[FFT.scala 34:12]
  wire [31:0] _GEN_841 = 11'h348 == cnt[10:0] ? $signed(32'sh474d) : $signed(_GEN_840); // @[FFT.scala 34:12]
  wire [31:0] _GEN_842 = 11'h349 == cnt[10:0] ? $signed(32'sh46ec) : $signed(_GEN_841); // @[FFT.scala 34:12]
  wire [31:0] _GEN_843 = 11'h34a == cnt[10:0] ? $signed(32'sh468c) : $signed(_GEN_842); // @[FFT.scala 34:12]
  wire [31:0] _GEN_844 = 11'h34b == cnt[10:0] ? $signed(32'sh462b) : $signed(_GEN_843); // @[FFT.scala 34:12]
  wire [31:0] _GEN_845 = 11'h34c == cnt[10:0] ? $signed(32'sh45cb) : $signed(_GEN_844); // @[FFT.scala 34:12]
  wire [31:0] _GEN_846 = 11'h34d == cnt[10:0] ? $signed(32'sh456a) : $signed(_GEN_845); // @[FFT.scala 34:12]
  wire [31:0] _GEN_847 = 11'h34e == cnt[10:0] ? $signed(32'sh4509) : $signed(_GEN_846); // @[FFT.scala 34:12]
  wire [31:0] _GEN_848 = 11'h34f == cnt[10:0] ? $signed(32'sh44a8) : $signed(_GEN_847); // @[FFT.scala 34:12]
  wire [31:0] _GEN_849 = 11'h350 == cnt[10:0] ? $signed(32'sh4447) : $signed(_GEN_848); // @[FFT.scala 34:12]
  wire [31:0] _GEN_850 = 11'h351 == cnt[10:0] ? $signed(32'sh43e6) : $signed(_GEN_849); // @[FFT.scala 34:12]
  wire [31:0] _GEN_851 = 11'h352 == cnt[10:0] ? $signed(32'sh4385) : $signed(_GEN_850); // @[FFT.scala 34:12]
  wire [31:0] _GEN_852 = 11'h353 == cnt[10:0] ? $signed(32'sh4324) : $signed(_GEN_851); // @[FFT.scala 34:12]
  wire [31:0] _GEN_853 = 11'h354 == cnt[10:0] ? $signed(32'sh42c3) : $signed(_GEN_852); // @[FFT.scala 34:12]
  wire [31:0] _GEN_854 = 11'h355 == cnt[10:0] ? $signed(32'sh4262) : $signed(_GEN_853); // @[FFT.scala 34:12]
  wire [31:0] _GEN_855 = 11'h356 == cnt[10:0] ? $signed(32'sh4201) : $signed(_GEN_854); // @[FFT.scala 34:12]
  wire [31:0] _GEN_856 = 11'h357 == cnt[10:0] ? $signed(32'sh41a0) : $signed(_GEN_855); // @[FFT.scala 34:12]
  wire [31:0] _GEN_857 = 11'h358 == cnt[10:0] ? $signed(32'sh413f) : $signed(_GEN_856); // @[FFT.scala 34:12]
  wire [31:0] _GEN_858 = 11'h359 == cnt[10:0] ? $signed(32'sh40de) : $signed(_GEN_857); // @[FFT.scala 34:12]
  wire [31:0] _GEN_859 = 11'h35a == cnt[10:0] ? $signed(32'sh407c) : $signed(_GEN_858); // @[FFT.scala 34:12]
  wire [31:0] _GEN_860 = 11'h35b == cnt[10:0] ? $signed(32'sh401b) : $signed(_GEN_859); // @[FFT.scala 34:12]
  wire [31:0] _GEN_861 = 11'h35c == cnt[10:0] ? $signed(32'sh3fba) : $signed(_GEN_860); // @[FFT.scala 34:12]
  wire [31:0] _GEN_862 = 11'h35d == cnt[10:0] ? $signed(32'sh3f58) : $signed(_GEN_861); // @[FFT.scala 34:12]
  wire [31:0] _GEN_863 = 11'h35e == cnt[10:0] ? $signed(32'sh3ef7) : $signed(_GEN_862); // @[FFT.scala 34:12]
  wire [31:0] _GEN_864 = 11'h35f == cnt[10:0] ? $signed(32'sh3e95) : $signed(_GEN_863); // @[FFT.scala 34:12]
  wire [31:0] _GEN_865 = 11'h360 == cnt[10:0] ? $signed(32'sh3e34) : $signed(_GEN_864); // @[FFT.scala 34:12]
  wire [31:0] _GEN_866 = 11'h361 == cnt[10:0] ? $signed(32'sh3dd2) : $signed(_GEN_865); // @[FFT.scala 34:12]
  wire [31:0] _GEN_867 = 11'h362 == cnt[10:0] ? $signed(32'sh3d71) : $signed(_GEN_866); // @[FFT.scala 34:12]
  wire [31:0] _GEN_868 = 11'h363 == cnt[10:0] ? $signed(32'sh3d0f) : $signed(_GEN_867); // @[FFT.scala 34:12]
  wire [31:0] _GEN_869 = 11'h364 == cnt[10:0] ? $signed(32'sh3cae) : $signed(_GEN_868); // @[FFT.scala 34:12]
  wire [31:0] _GEN_870 = 11'h365 == cnt[10:0] ? $signed(32'sh3c4c) : $signed(_GEN_869); // @[FFT.scala 34:12]
  wire [31:0] _GEN_871 = 11'h366 == cnt[10:0] ? $signed(32'sh3bea) : $signed(_GEN_870); // @[FFT.scala 34:12]
  wire [31:0] _GEN_872 = 11'h367 == cnt[10:0] ? $signed(32'sh3b88) : $signed(_GEN_871); // @[FFT.scala 34:12]
  wire [31:0] _GEN_873 = 11'h368 == cnt[10:0] ? $signed(32'sh3b27) : $signed(_GEN_872); // @[FFT.scala 34:12]
  wire [31:0] _GEN_874 = 11'h369 == cnt[10:0] ? $signed(32'sh3ac5) : $signed(_GEN_873); // @[FFT.scala 34:12]
  wire [31:0] _GEN_875 = 11'h36a == cnt[10:0] ? $signed(32'sh3a63) : $signed(_GEN_874); // @[FFT.scala 34:12]
  wire [31:0] _GEN_876 = 11'h36b == cnt[10:0] ? $signed(32'sh3a01) : $signed(_GEN_875); // @[FFT.scala 34:12]
  wire [31:0] _GEN_877 = 11'h36c == cnt[10:0] ? $signed(32'sh399f) : $signed(_GEN_876); // @[FFT.scala 34:12]
  wire [31:0] _GEN_878 = 11'h36d == cnt[10:0] ? $signed(32'sh393d) : $signed(_GEN_877); // @[FFT.scala 34:12]
  wire [31:0] _GEN_879 = 11'h36e == cnt[10:0] ? $signed(32'sh38db) : $signed(_GEN_878); // @[FFT.scala 34:12]
  wire [31:0] _GEN_880 = 11'h36f == cnt[10:0] ? $signed(32'sh3879) : $signed(_GEN_879); // @[FFT.scala 34:12]
  wire [31:0] _GEN_881 = 11'h370 == cnt[10:0] ? $signed(32'sh3817) : $signed(_GEN_880); // @[FFT.scala 34:12]
  wire [31:0] _GEN_882 = 11'h371 == cnt[10:0] ? $signed(32'sh37b5) : $signed(_GEN_881); // @[FFT.scala 34:12]
  wire [31:0] _GEN_883 = 11'h372 == cnt[10:0] ? $signed(32'sh3753) : $signed(_GEN_882); // @[FFT.scala 34:12]
  wire [31:0] _GEN_884 = 11'h373 == cnt[10:0] ? $signed(32'sh36f1) : $signed(_GEN_883); // @[FFT.scala 34:12]
  wire [31:0] _GEN_885 = 11'h374 == cnt[10:0] ? $signed(32'sh368e) : $signed(_GEN_884); // @[FFT.scala 34:12]
  wire [31:0] _GEN_886 = 11'h375 == cnt[10:0] ? $signed(32'sh362c) : $signed(_GEN_885); // @[FFT.scala 34:12]
  wire [31:0] _GEN_887 = 11'h376 == cnt[10:0] ? $signed(32'sh35ca) : $signed(_GEN_886); // @[FFT.scala 34:12]
  wire [31:0] _GEN_888 = 11'h377 == cnt[10:0] ? $signed(32'sh3568) : $signed(_GEN_887); // @[FFT.scala 34:12]
  wire [31:0] _GEN_889 = 11'h378 == cnt[10:0] ? $signed(32'sh3505) : $signed(_GEN_888); // @[FFT.scala 34:12]
  wire [31:0] _GEN_890 = 11'h379 == cnt[10:0] ? $signed(32'sh34a3) : $signed(_GEN_889); // @[FFT.scala 34:12]
  wire [31:0] _GEN_891 = 11'h37a == cnt[10:0] ? $signed(32'sh3440) : $signed(_GEN_890); // @[FFT.scala 34:12]
  wire [31:0] _GEN_892 = 11'h37b == cnt[10:0] ? $signed(32'sh33de) : $signed(_GEN_891); // @[FFT.scala 34:12]
  wire [31:0] _GEN_893 = 11'h37c == cnt[10:0] ? $signed(32'sh337c) : $signed(_GEN_892); // @[FFT.scala 34:12]
  wire [31:0] _GEN_894 = 11'h37d == cnt[10:0] ? $signed(32'sh3319) : $signed(_GEN_893); // @[FFT.scala 34:12]
  wire [31:0] _GEN_895 = 11'h37e == cnt[10:0] ? $signed(32'sh32b7) : $signed(_GEN_894); // @[FFT.scala 34:12]
  wire [31:0] _GEN_896 = 11'h37f == cnt[10:0] ? $signed(32'sh3254) : $signed(_GEN_895); // @[FFT.scala 34:12]
  wire [31:0] _GEN_897 = 11'h380 == cnt[10:0] ? $signed(32'sh31f1) : $signed(_GEN_896); // @[FFT.scala 34:12]
  wire [31:0] _GEN_898 = 11'h381 == cnt[10:0] ? $signed(32'sh318f) : $signed(_GEN_897); // @[FFT.scala 34:12]
  wire [31:0] _GEN_899 = 11'h382 == cnt[10:0] ? $signed(32'sh312c) : $signed(_GEN_898); // @[FFT.scala 34:12]
  wire [31:0] _GEN_900 = 11'h383 == cnt[10:0] ? $signed(32'sh30ca) : $signed(_GEN_899); // @[FFT.scala 34:12]
  wire [31:0] _GEN_901 = 11'h384 == cnt[10:0] ? $signed(32'sh3067) : $signed(_GEN_900); // @[FFT.scala 34:12]
  wire [31:0] _GEN_902 = 11'h385 == cnt[10:0] ? $signed(32'sh3004) : $signed(_GEN_901); // @[FFT.scala 34:12]
  wire [31:0] _GEN_903 = 11'h386 == cnt[10:0] ? $signed(32'sh2fa1) : $signed(_GEN_902); // @[FFT.scala 34:12]
  wire [31:0] _GEN_904 = 11'h387 == cnt[10:0] ? $signed(32'sh2f3f) : $signed(_GEN_903); // @[FFT.scala 34:12]
  wire [31:0] _GEN_905 = 11'h388 == cnt[10:0] ? $signed(32'sh2edc) : $signed(_GEN_904); // @[FFT.scala 34:12]
  wire [31:0] _GEN_906 = 11'h389 == cnt[10:0] ? $signed(32'sh2e79) : $signed(_GEN_905); // @[FFT.scala 34:12]
  wire [31:0] _GEN_907 = 11'h38a == cnt[10:0] ? $signed(32'sh2e16) : $signed(_GEN_906); // @[FFT.scala 34:12]
  wire [31:0] _GEN_908 = 11'h38b == cnt[10:0] ? $signed(32'sh2db3) : $signed(_GEN_907); // @[FFT.scala 34:12]
  wire [31:0] _GEN_909 = 11'h38c == cnt[10:0] ? $signed(32'sh2d50) : $signed(_GEN_908); // @[FFT.scala 34:12]
  wire [31:0] _GEN_910 = 11'h38d == cnt[10:0] ? $signed(32'sh2ced) : $signed(_GEN_909); // @[FFT.scala 34:12]
  wire [31:0] _GEN_911 = 11'h38e == cnt[10:0] ? $signed(32'sh2c8a) : $signed(_GEN_910); // @[FFT.scala 34:12]
  wire [31:0] _GEN_912 = 11'h38f == cnt[10:0] ? $signed(32'sh2c27) : $signed(_GEN_911); // @[FFT.scala 34:12]
  wire [31:0] _GEN_913 = 11'h390 == cnt[10:0] ? $signed(32'sh2bc4) : $signed(_GEN_912); // @[FFT.scala 34:12]
  wire [31:0] _GEN_914 = 11'h391 == cnt[10:0] ? $signed(32'sh2b61) : $signed(_GEN_913); // @[FFT.scala 34:12]
  wire [31:0] _GEN_915 = 11'h392 == cnt[10:0] ? $signed(32'sh2afe) : $signed(_GEN_914); // @[FFT.scala 34:12]
  wire [31:0] _GEN_916 = 11'h393 == cnt[10:0] ? $signed(32'sh2a9b) : $signed(_GEN_915); // @[FFT.scala 34:12]
  wire [31:0] _GEN_917 = 11'h394 == cnt[10:0] ? $signed(32'sh2a38) : $signed(_GEN_916); // @[FFT.scala 34:12]
  wire [31:0] _GEN_918 = 11'h395 == cnt[10:0] ? $signed(32'sh29d5) : $signed(_GEN_917); // @[FFT.scala 34:12]
  wire [31:0] _GEN_919 = 11'h396 == cnt[10:0] ? $signed(32'sh2971) : $signed(_GEN_918); // @[FFT.scala 34:12]
  wire [31:0] _GEN_920 = 11'h397 == cnt[10:0] ? $signed(32'sh290e) : $signed(_GEN_919); // @[FFT.scala 34:12]
  wire [31:0] _GEN_921 = 11'h398 == cnt[10:0] ? $signed(32'sh28ab) : $signed(_GEN_920); // @[FFT.scala 34:12]
  wire [31:0] _GEN_922 = 11'h399 == cnt[10:0] ? $signed(32'sh2848) : $signed(_GEN_921); // @[FFT.scala 34:12]
  wire [31:0] _GEN_923 = 11'h39a == cnt[10:0] ? $signed(32'sh27e4) : $signed(_GEN_922); // @[FFT.scala 34:12]
  wire [31:0] _GEN_924 = 11'h39b == cnt[10:0] ? $signed(32'sh2781) : $signed(_GEN_923); // @[FFT.scala 34:12]
  wire [31:0] _GEN_925 = 11'h39c == cnt[10:0] ? $signed(32'sh271e) : $signed(_GEN_924); // @[FFT.scala 34:12]
  wire [31:0] _GEN_926 = 11'h39d == cnt[10:0] ? $signed(32'sh26ba) : $signed(_GEN_925); // @[FFT.scala 34:12]
  wire [31:0] _GEN_927 = 11'h39e == cnt[10:0] ? $signed(32'sh2657) : $signed(_GEN_926); // @[FFT.scala 34:12]
  wire [31:0] _GEN_928 = 11'h39f == cnt[10:0] ? $signed(32'sh25f4) : $signed(_GEN_927); // @[FFT.scala 34:12]
  wire [31:0] _GEN_929 = 11'h3a0 == cnt[10:0] ? $signed(32'sh2590) : $signed(_GEN_928); // @[FFT.scala 34:12]
  wire [31:0] _GEN_930 = 11'h3a1 == cnt[10:0] ? $signed(32'sh252d) : $signed(_GEN_929); // @[FFT.scala 34:12]
  wire [31:0] _GEN_931 = 11'h3a2 == cnt[10:0] ? $signed(32'sh24c9) : $signed(_GEN_930); // @[FFT.scala 34:12]
  wire [31:0] _GEN_932 = 11'h3a3 == cnt[10:0] ? $signed(32'sh2466) : $signed(_GEN_931); // @[FFT.scala 34:12]
  wire [31:0] _GEN_933 = 11'h3a4 == cnt[10:0] ? $signed(32'sh2402) : $signed(_GEN_932); // @[FFT.scala 34:12]
  wire [31:0] _GEN_934 = 11'h3a5 == cnt[10:0] ? $signed(32'sh239f) : $signed(_GEN_933); // @[FFT.scala 34:12]
  wire [31:0] _GEN_935 = 11'h3a6 == cnt[10:0] ? $signed(32'sh233b) : $signed(_GEN_934); // @[FFT.scala 34:12]
  wire [31:0] _GEN_936 = 11'h3a7 == cnt[10:0] ? $signed(32'sh22d7) : $signed(_GEN_935); // @[FFT.scala 34:12]
  wire [31:0] _GEN_937 = 11'h3a8 == cnt[10:0] ? $signed(32'sh2274) : $signed(_GEN_936); // @[FFT.scala 34:12]
  wire [31:0] _GEN_938 = 11'h3a9 == cnt[10:0] ? $signed(32'sh2210) : $signed(_GEN_937); // @[FFT.scala 34:12]
  wire [31:0] _GEN_939 = 11'h3aa == cnt[10:0] ? $signed(32'sh21ad) : $signed(_GEN_938); // @[FFT.scala 34:12]
  wire [31:0] _GEN_940 = 11'h3ab == cnt[10:0] ? $signed(32'sh2149) : $signed(_GEN_939); // @[FFT.scala 34:12]
  wire [31:0] _GEN_941 = 11'h3ac == cnt[10:0] ? $signed(32'sh20e5) : $signed(_GEN_940); // @[FFT.scala 34:12]
  wire [31:0] _GEN_942 = 11'h3ad == cnt[10:0] ? $signed(32'sh2082) : $signed(_GEN_941); // @[FFT.scala 34:12]
  wire [31:0] _GEN_943 = 11'h3ae == cnt[10:0] ? $signed(32'sh201e) : $signed(_GEN_942); // @[FFT.scala 34:12]
  wire [31:0] _GEN_944 = 11'h3af == cnt[10:0] ? $signed(32'sh1fba) : $signed(_GEN_943); // @[FFT.scala 34:12]
  wire [31:0] _GEN_945 = 11'h3b0 == cnt[10:0] ? $signed(32'sh1f56) : $signed(_GEN_944); // @[FFT.scala 34:12]
  wire [31:0] _GEN_946 = 11'h3b1 == cnt[10:0] ? $signed(32'sh1ef3) : $signed(_GEN_945); // @[FFT.scala 34:12]
  wire [31:0] _GEN_947 = 11'h3b2 == cnt[10:0] ? $signed(32'sh1e8f) : $signed(_GEN_946); // @[FFT.scala 34:12]
  wire [31:0] _GEN_948 = 11'h3b3 == cnt[10:0] ? $signed(32'sh1e2b) : $signed(_GEN_947); // @[FFT.scala 34:12]
  wire [31:0] _GEN_949 = 11'h3b4 == cnt[10:0] ? $signed(32'sh1dc7) : $signed(_GEN_948); // @[FFT.scala 34:12]
  wire [31:0] _GEN_950 = 11'h3b5 == cnt[10:0] ? $signed(32'sh1d63) : $signed(_GEN_949); // @[FFT.scala 34:12]
  wire [31:0] _GEN_951 = 11'h3b6 == cnt[10:0] ? $signed(32'sh1cff) : $signed(_GEN_950); // @[FFT.scala 34:12]
  wire [31:0] _GEN_952 = 11'h3b7 == cnt[10:0] ? $signed(32'sh1c9b) : $signed(_GEN_951); // @[FFT.scala 34:12]
  wire [31:0] _GEN_953 = 11'h3b8 == cnt[10:0] ? $signed(32'sh1c38) : $signed(_GEN_952); // @[FFT.scala 34:12]
  wire [31:0] _GEN_954 = 11'h3b9 == cnt[10:0] ? $signed(32'sh1bd4) : $signed(_GEN_953); // @[FFT.scala 34:12]
  wire [31:0] _GEN_955 = 11'h3ba == cnt[10:0] ? $signed(32'sh1b70) : $signed(_GEN_954); // @[FFT.scala 34:12]
  wire [31:0] _GEN_956 = 11'h3bb == cnt[10:0] ? $signed(32'sh1b0c) : $signed(_GEN_955); // @[FFT.scala 34:12]
  wire [31:0] _GEN_957 = 11'h3bc == cnt[10:0] ? $signed(32'sh1aa8) : $signed(_GEN_956); // @[FFT.scala 34:12]
  wire [31:0] _GEN_958 = 11'h3bd == cnt[10:0] ? $signed(32'sh1a44) : $signed(_GEN_957); // @[FFT.scala 34:12]
  wire [31:0] _GEN_959 = 11'h3be == cnt[10:0] ? $signed(32'sh19e0) : $signed(_GEN_958); // @[FFT.scala 34:12]
  wire [31:0] _GEN_960 = 11'h3bf == cnt[10:0] ? $signed(32'sh197c) : $signed(_GEN_959); // @[FFT.scala 34:12]
  wire [31:0] _GEN_961 = 11'h3c0 == cnt[10:0] ? $signed(32'sh1918) : $signed(_GEN_960); // @[FFT.scala 34:12]
  wire [31:0] _GEN_962 = 11'h3c1 == cnt[10:0] ? $signed(32'sh18b4) : $signed(_GEN_961); // @[FFT.scala 34:12]
  wire [31:0] _GEN_963 = 11'h3c2 == cnt[10:0] ? $signed(32'sh1850) : $signed(_GEN_962); // @[FFT.scala 34:12]
  wire [31:0] _GEN_964 = 11'h3c3 == cnt[10:0] ? $signed(32'sh17eb) : $signed(_GEN_963); // @[FFT.scala 34:12]
  wire [31:0] _GEN_965 = 11'h3c4 == cnt[10:0] ? $signed(32'sh1787) : $signed(_GEN_964); // @[FFT.scala 34:12]
  wire [31:0] _GEN_966 = 11'h3c5 == cnt[10:0] ? $signed(32'sh1723) : $signed(_GEN_965); // @[FFT.scala 34:12]
  wire [31:0] _GEN_967 = 11'h3c6 == cnt[10:0] ? $signed(32'sh16bf) : $signed(_GEN_966); // @[FFT.scala 34:12]
  wire [31:0] _GEN_968 = 11'h3c7 == cnt[10:0] ? $signed(32'sh165b) : $signed(_GEN_967); // @[FFT.scala 34:12]
  wire [31:0] _GEN_969 = 11'h3c8 == cnt[10:0] ? $signed(32'sh15f7) : $signed(_GEN_968); // @[FFT.scala 34:12]
  wire [31:0] _GEN_970 = 11'h3c9 == cnt[10:0] ? $signed(32'sh1593) : $signed(_GEN_969); // @[FFT.scala 34:12]
  wire [31:0] _GEN_971 = 11'h3ca == cnt[10:0] ? $signed(32'sh152e) : $signed(_GEN_970); // @[FFT.scala 34:12]
  wire [31:0] _GEN_972 = 11'h3cb == cnt[10:0] ? $signed(32'sh14ca) : $signed(_GEN_971); // @[FFT.scala 34:12]
  wire [31:0] _GEN_973 = 11'h3cc == cnt[10:0] ? $signed(32'sh1466) : $signed(_GEN_972); // @[FFT.scala 34:12]
  wire [31:0] _GEN_974 = 11'h3cd == cnt[10:0] ? $signed(32'sh1402) : $signed(_GEN_973); // @[FFT.scala 34:12]
  wire [31:0] _GEN_975 = 11'h3ce == cnt[10:0] ? $signed(32'sh139e) : $signed(_GEN_974); // @[FFT.scala 34:12]
  wire [31:0] _GEN_976 = 11'h3cf == cnt[10:0] ? $signed(32'sh1339) : $signed(_GEN_975); // @[FFT.scala 34:12]
  wire [31:0] _GEN_977 = 11'h3d0 == cnt[10:0] ? $signed(32'sh12d5) : $signed(_GEN_976); // @[FFT.scala 34:12]
  wire [31:0] _GEN_978 = 11'h3d1 == cnt[10:0] ? $signed(32'sh1271) : $signed(_GEN_977); // @[FFT.scala 34:12]
  wire [31:0] _GEN_979 = 11'h3d2 == cnt[10:0] ? $signed(32'sh120d) : $signed(_GEN_978); // @[FFT.scala 34:12]
  wire [31:0] _GEN_980 = 11'h3d3 == cnt[10:0] ? $signed(32'sh11a8) : $signed(_GEN_979); // @[FFT.scala 34:12]
  wire [31:0] _GEN_981 = 11'h3d4 == cnt[10:0] ? $signed(32'sh1144) : $signed(_GEN_980); // @[FFT.scala 34:12]
  wire [31:0] _GEN_982 = 11'h3d5 == cnt[10:0] ? $signed(32'sh10e0) : $signed(_GEN_981); // @[FFT.scala 34:12]
  wire [31:0] _GEN_983 = 11'h3d6 == cnt[10:0] ? $signed(32'sh107b) : $signed(_GEN_982); // @[FFT.scala 34:12]
  wire [31:0] _GEN_984 = 11'h3d7 == cnt[10:0] ? $signed(32'sh1017) : $signed(_GEN_983); // @[FFT.scala 34:12]
  wire [31:0] _GEN_985 = 11'h3d8 == cnt[10:0] ? $signed(32'shfb3) : $signed(_GEN_984); // @[FFT.scala 34:12]
  wire [31:0] _GEN_986 = 11'h3d9 == cnt[10:0] ? $signed(32'shf4e) : $signed(_GEN_985); // @[FFT.scala 34:12]
  wire [31:0] _GEN_987 = 11'h3da == cnt[10:0] ? $signed(32'sheea) : $signed(_GEN_986); // @[FFT.scala 34:12]
  wire [31:0] _GEN_988 = 11'h3db == cnt[10:0] ? $signed(32'she86) : $signed(_GEN_987); // @[FFT.scala 34:12]
  wire [31:0] _GEN_989 = 11'h3dc == cnt[10:0] ? $signed(32'she21) : $signed(_GEN_988); // @[FFT.scala 34:12]
  wire [31:0] _GEN_990 = 11'h3dd == cnt[10:0] ? $signed(32'shdbd) : $signed(_GEN_989); // @[FFT.scala 34:12]
  wire [31:0] _GEN_991 = 11'h3de == cnt[10:0] ? $signed(32'shd59) : $signed(_GEN_990); // @[FFT.scala 34:12]
  wire [31:0] _GEN_992 = 11'h3df == cnt[10:0] ? $signed(32'shcf4) : $signed(_GEN_991); // @[FFT.scala 34:12]
  wire [31:0] _GEN_993 = 11'h3e0 == cnt[10:0] ? $signed(32'shc90) : $signed(_GEN_992); // @[FFT.scala 34:12]
  wire [31:0] _GEN_994 = 11'h3e1 == cnt[10:0] ? $signed(32'shc2b) : $signed(_GEN_993); // @[FFT.scala 34:12]
  wire [31:0] _GEN_995 = 11'h3e2 == cnt[10:0] ? $signed(32'shbc7) : $signed(_GEN_994); // @[FFT.scala 34:12]
  wire [31:0] _GEN_996 = 11'h3e3 == cnt[10:0] ? $signed(32'shb62) : $signed(_GEN_995); // @[FFT.scala 34:12]
  wire [31:0] _GEN_997 = 11'h3e4 == cnt[10:0] ? $signed(32'shafe) : $signed(_GEN_996); // @[FFT.scala 34:12]
  wire [31:0] _GEN_998 = 11'h3e5 == cnt[10:0] ? $signed(32'sha9a) : $signed(_GEN_997); // @[FFT.scala 34:12]
  wire [31:0] _GEN_999 = 11'h3e6 == cnt[10:0] ? $signed(32'sha35) : $signed(_GEN_998); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1000 = 11'h3e7 == cnt[10:0] ? $signed(32'sh9d1) : $signed(_GEN_999); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1001 = 11'h3e8 == cnt[10:0] ? $signed(32'sh96c) : $signed(_GEN_1000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1002 = 11'h3e9 == cnt[10:0] ? $signed(32'sh908) : $signed(_GEN_1001); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1003 = 11'h3ea == cnt[10:0] ? $signed(32'sh8a3) : $signed(_GEN_1002); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1004 = 11'h3eb == cnt[10:0] ? $signed(32'sh83f) : $signed(_GEN_1003); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1005 = 11'h3ec == cnt[10:0] ? $signed(32'sh7da) : $signed(_GEN_1004); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1006 = 11'h3ed == cnt[10:0] ? $signed(32'sh776) : $signed(_GEN_1005); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1007 = 11'h3ee == cnt[10:0] ? $signed(32'sh711) : $signed(_GEN_1006); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1008 = 11'h3ef == cnt[10:0] ? $signed(32'sh6ad) : $signed(_GEN_1007); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1009 = 11'h3f0 == cnt[10:0] ? $signed(32'sh648) : $signed(_GEN_1008); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1010 = 11'h3f1 == cnt[10:0] ? $signed(32'sh5e4) : $signed(_GEN_1009); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1011 = 11'h3f2 == cnt[10:0] ? $signed(32'sh57f) : $signed(_GEN_1010); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1012 = 11'h3f3 == cnt[10:0] ? $signed(32'sh51b) : $signed(_GEN_1011); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1013 = 11'h3f4 == cnt[10:0] ? $signed(32'sh4b6) : $signed(_GEN_1012); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1014 = 11'h3f5 == cnt[10:0] ? $signed(32'sh452) : $signed(_GEN_1013); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1015 = 11'h3f6 == cnt[10:0] ? $signed(32'sh3ed) : $signed(_GEN_1014); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1016 = 11'h3f7 == cnt[10:0] ? $signed(32'sh389) : $signed(_GEN_1015); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1017 = 11'h3f8 == cnt[10:0] ? $signed(32'sh324) : $signed(_GEN_1016); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1018 = 11'h3f9 == cnt[10:0] ? $signed(32'sh2c0) : $signed(_GEN_1017); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1019 = 11'h3fa == cnt[10:0] ? $signed(32'sh25b) : $signed(_GEN_1018); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1020 = 11'h3fb == cnt[10:0] ? $signed(32'sh1f7) : $signed(_GEN_1019); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1021 = 11'h3fc == cnt[10:0] ? $signed(32'sh192) : $signed(_GEN_1020); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1022 = 11'h3fd == cnt[10:0] ? $signed(32'sh12e) : $signed(_GEN_1021); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1023 = 11'h3fe == cnt[10:0] ? $signed(32'shc9) : $signed(_GEN_1022); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1024 = 11'h3ff == cnt[10:0] ? $signed(32'sh65) : $signed(_GEN_1023); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1025 = 11'h400 == cnt[10:0] ? $signed(32'sh0) : $signed(_GEN_1024); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1026 = 11'h401 == cnt[10:0] ? $signed(-32'sh65) : $signed(_GEN_1025); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1027 = 11'h402 == cnt[10:0] ? $signed(-32'shc9) : $signed(_GEN_1026); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1028 = 11'h403 == cnt[10:0] ? $signed(-32'sh12e) : $signed(_GEN_1027); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1029 = 11'h404 == cnt[10:0] ? $signed(-32'sh192) : $signed(_GEN_1028); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1030 = 11'h405 == cnt[10:0] ? $signed(-32'sh1f7) : $signed(_GEN_1029); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1031 = 11'h406 == cnt[10:0] ? $signed(-32'sh25b) : $signed(_GEN_1030); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1032 = 11'h407 == cnt[10:0] ? $signed(-32'sh2c0) : $signed(_GEN_1031); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1033 = 11'h408 == cnt[10:0] ? $signed(-32'sh324) : $signed(_GEN_1032); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1034 = 11'h409 == cnt[10:0] ? $signed(-32'sh389) : $signed(_GEN_1033); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1035 = 11'h40a == cnt[10:0] ? $signed(-32'sh3ed) : $signed(_GEN_1034); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1036 = 11'h40b == cnt[10:0] ? $signed(-32'sh452) : $signed(_GEN_1035); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1037 = 11'h40c == cnt[10:0] ? $signed(-32'sh4b6) : $signed(_GEN_1036); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1038 = 11'h40d == cnt[10:0] ? $signed(-32'sh51b) : $signed(_GEN_1037); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1039 = 11'h40e == cnt[10:0] ? $signed(-32'sh57f) : $signed(_GEN_1038); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1040 = 11'h40f == cnt[10:0] ? $signed(-32'sh5e4) : $signed(_GEN_1039); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1041 = 11'h410 == cnt[10:0] ? $signed(-32'sh648) : $signed(_GEN_1040); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1042 = 11'h411 == cnt[10:0] ? $signed(-32'sh6ad) : $signed(_GEN_1041); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1043 = 11'h412 == cnt[10:0] ? $signed(-32'sh711) : $signed(_GEN_1042); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1044 = 11'h413 == cnt[10:0] ? $signed(-32'sh776) : $signed(_GEN_1043); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1045 = 11'h414 == cnt[10:0] ? $signed(-32'sh7da) : $signed(_GEN_1044); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1046 = 11'h415 == cnt[10:0] ? $signed(-32'sh83f) : $signed(_GEN_1045); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1047 = 11'h416 == cnt[10:0] ? $signed(-32'sh8a3) : $signed(_GEN_1046); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1048 = 11'h417 == cnt[10:0] ? $signed(-32'sh908) : $signed(_GEN_1047); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1049 = 11'h418 == cnt[10:0] ? $signed(-32'sh96c) : $signed(_GEN_1048); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1050 = 11'h419 == cnt[10:0] ? $signed(-32'sh9d1) : $signed(_GEN_1049); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1051 = 11'h41a == cnt[10:0] ? $signed(-32'sha35) : $signed(_GEN_1050); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1052 = 11'h41b == cnt[10:0] ? $signed(-32'sha9a) : $signed(_GEN_1051); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1053 = 11'h41c == cnt[10:0] ? $signed(-32'shafe) : $signed(_GEN_1052); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1054 = 11'h41d == cnt[10:0] ? $signed(-32'shb62) : $signed(_GEN_1053); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1055 = 11'h41e == cnt[10:0] ? $signed(-32'shbc7) : $signed(_GEN_1054); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1056 = 11'h41f == cnt[10:0] ? $signed(-32'shc2b) : $signed(_GEN_1055); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1057 = 11'h420 == cnt[10:0] ? $signed(-32'shc90) : $signed(_GEN_1056); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1058 = 11'h421 == cnt[10:0] ? $signed(-32'shcf4) : $signed(_GEN_1057); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1059 = 11'h422 == cnt[10:0] ? $signed(-32'shd59) : $signed(_GEN_1058); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1060 = 11'h423 == cnt[10:0] ? $signed(-32'shdbd) : $signed(_GEN_1059); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1061 = 11'h424 == cnt[10:0] ? $signed(-32'she21) : $signed(_GEN_1060); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1062 = 11'h425 == cnt[10:0] ? $signed(-32'she86) : $signed(_GEN_1061); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1063 = 11'h426 == cnt[10:0] ? $signed(-32'sheea) : $signed(_GEN_1062); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1064 = 11'h427 == cnt[10:0] ? $signed(-32'shf4e) : $signed(_GEN_1063); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1065 = 11'h428 == cnt[10:0] ? $signed(-32'shfb3) : $signed(_GEN_1064); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1066 = 11'h429 == cnt[10:0] ? $signed(-32'sh1017) : $signed(_GEN_1065); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1067 = 11'h42a == cnt[10:0] ? $signed(-32'sh107b) : $signed(_GEN_1066); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1068 = 11'h42b == cnt[10:0] ? $signed(-32'sh10e0) : $signed(_GEN_1067); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1069 = 11'h42c == cnt[10:0] ? $signed(-32'sh1144) : $signed(_GEN_1068); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1070 = 11'h42d == cnt[10:0] ? $signed(-32'sh11a8) : $signed(_GEN_1069); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1071 = 11'h42e == cnt[10:0] ? $signed(-32'sh120d) : $signed(_GEN_1070); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1072 = 11'h42f == cnt[10:0] ? $signed(-32'sh1271) : $signed(_GEN_1071); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1073 = 11'h430 == cnt[10:0] ? $signed(-32'sh12d5) : $signed(_GEN_1072); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1074 = 11'h431 == cnt[10:0] ? $signed(-32'sh1339) : $signed(_GEN_1073); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1075 = 11'h432 == cnt[10:0] ? $signed(-32'sh139e) : $signed(_GEN_1074); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1076 = 11'h433 == cnt[10:0] ? $signed(-32'sh1402) : $signed(_GEN_1075); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1077 = 11'h434 == cnt[10:0] ? $signed(-32'sh1466) : $signed(_GEN_1076); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1078 = 11'h435 == cnt[10:0] ? $signed(-32'sh14ca) : $signed(_GEN_1077); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1079 = 11'h436 == cnt[10:0] ? $signed(-32'sh152e) : $signed(_GEN_1078); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1080 = 11'h437 == cnt[10:0] ? $signed(-32'sh1593) : $signed(_GEN_1079); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1081 = 11'h438 == cnt[10:0] ? $signed(-32'sh15f7) : $signed(_GEN_1080); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1082 = 11'h439 == cnt[10:0] ? $signed(-32'sh165b) : $signed(_GEN_1081); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1083 = 11'h43a == cnt[10:0] ? $signed(-32'sh16bf) : $signed(_GEN_1082); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1084 = 11'h43b == cnt[10:0] ? $signed(-32'sh1723) : $signed(_GEN_1083); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1085 = 11'h43c == cnt[10:0] ? $signed(-32'sh1787) : $signed(_GEN_1084); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1086 = 11'h43d == cnt[10:0] ? $signed(-32'sh17eb) : $signed(_GEN_1085); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1087 = 11'h43e == cnt[10:0] ? $signed(-32'sh1850) : $signed(_GEN_1086); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1088 = 11'h43f == cnt[10:0] ? $signed(-32'sh18b4) : $signed(_GEN_1087); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1089 = 11'h440 == cnt[10:0] ? $signed(-32'sh1918) : $signed(_GEN_1088); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1090 = 11'h441 == cnt[10:0] ? $signed(-32'sh197c) : $signed(_GEN_1089); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1091 = 11'h442 == cnt[10:0] ? $signed(-32'sh19e0) : $signed(_GEN_1090); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1092 = 11'h443 == cnt[10:0] ? $signed(-32'sh1a44) : $signed(_GEN_1091); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1093 = 11'h444 == cnt[10:0] ? $signed(-32'sh1aa8) : $signed(_GEN_1092); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1094 = 11'h445 == cnt[10:0] ? $signed(-32'sh1b0c) : $signed(_GEN_1093); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1095 = 11'h446 == cnt[10:0] ? $signed(-32'sh1b70) : $signed(_GEN_1094); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1096 = 11'h447 == cnt[10:0] ? $signed(-32'sh1bd4) : $signed(_GEN_1095); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1097 = 11'h448 == cnt[10:0] ? $signed(-32'sh1c38) : $signed(_GEN_1096); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1098 = 11'h449 == cnt[10:0] ? $signed(-32'sh1c9b) : $signed(_GEN_1097); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1099 = 11'h44a == cnt[10:0] ? $signed(-32'sh1cff) : $signed(_GEN_1098); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1100 = 11'h44b == cnt[10:0] ? $signed(-32'sh1d63) : $signed(_GEN_1099); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1101 = 11'h44c == cnt[10:0] ? $signed(-32'sh1dc7) : $signed(_GEN_1100); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1102 = 11'h44d == cnt[10:0] ? $signed(-32'sh1e2b) : $signed(_GEN_1101); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1103 = 11'h44e == cnt[10:0] ? $signed(-32'sh1e8f) : $signed(_GEN_1102); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1104 = 11'h44f == cnt[10:0] ? $signed(-32'sh1ef3) : $signed(_GEN_1103); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1105 = 11'h450 == cnt[10:0] ? $signed(-32'sh1f56) : $signed(_GEN_1104); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1106 = 11'h451 == cnt[10:0] ? $signed(-32'sh1fba) : $signed(_GEN_1105); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1107 = 11'h452 == cnt[10:0] ? $signed(-32'sh201e) : $signed(_GEN_1106); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1108 = 11'h453 == cnt[10:0] ? $signed(-32'sh2082) : $signed(_GEN_1107); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1109 = 11'h454 == cnt[10:0] ? $signed(-32'sh20e5) : $signed(_GEN_1108); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1110 = 11'h455 == cnt[10:0] ? $signed(-32'sh2149) : $signed(_GEN_1109); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1111 = 11'h456 == cnt[10:0] ? $signed(-32'sh21ad) : $signed(_GEN_1110); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1112 = 11'h457 == cnt[10:0] ? $signed(-32'sh2210) : $signed(_GEN_1111); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1113 = 11'h458 == cnt[10:0] ? $signed(-32'sh2274) : $signed(_GEN_1112); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1114 = 11'h459 == cnt[10:0] ? $signed(-32'sh22d7) : $signed(_GEN_1113); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1115 = 11'h45a == cnt[10:0] ? $signed(-32'sh233b) : $signed(_GEN_1114); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1116 = 11'h45b == cnt[10:0] ? $signed(-32'sh239f) : $signed(_GEN_1115); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1117 = 11'h45c == cnt[10:0] ? $signed(-32'sh2402) : $signed(_GEN_1116); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1118 = 11'h45d == cnt[10:0] ? $signed(-32'sh2466) : $signed(_GEN_1117); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1119 = 11'h45e == cnt[10:0] ? $signed(-32'sh24c9) : $signed(_GEN_1118); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1120 = 11'h45f == cnt[10:0] ? $signed(-32'sh252d) : $signed(_GEN_1119); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1121 = 11'h460 == cnt[10:0] ? $signed(-32'sh2590) : $signed(_GEN_1120); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1122 = 11'h461 == cnt[10:0] ? $signed(-32'sh25f4) : $signed(_GEN_1121); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1123 = 11'h462 == cnt[10:0] ? $signed(-32'sh2657) : $signed(_GEN_1122); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1124 = 11'h463 == cnt[10:0] ? $signed(-32'sh26ba) : $signed(_GEN_1123); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1125 = 11'h464 == cnt[10:0] ? $signed(-32'sh271e) : $signed(_GEN_1124); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1126 = 11'h465 == cnt[10:0] ? $signed(-32'sh2781) : $signed(_GEN_1125); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1127 = 11'h466 == cnt[10:0] ? $signed(-32'sh27e4) : $signed(_GEN_1126); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1128 = 11'h467 == cnt[10:0] ? $signed(-32'sh2848) : $signed(_GEN_1127); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1129 = 11'h468 == cnt[10:0] ? $signed(-32'sh28ab) : $signed(_GEN_1128); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1130 = 11'h469 == cnt[10:0] ? $signed(-32'sh290e) : $signed(_GEN_1129); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1131 = 11'h46a == cnt[10:0] ? $signed(-32'sh2971) : $signed(_GEN_1130); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1132 = 11'h46b == cnt[10:0] ? $signed(-32'sh29d5) : $signed(_GEN_1131); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1133 = 11'h46c == cnt[10:0] ? $signed(-32'sh2a38) : $signed(_GEN_1132); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1134 = 11'h46d == cnt[10:0] ? $signed(-32'sh2a9b) : $signed(_GEN_1133); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1135 = 11'h46e == cnt[10:0] ? $signed(-32'sh2afe) : $signed(_GEN_1134); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1136 = 11'h46f == cnt[10:0] ? $signed(-32'sh2b61) : $signed(_GEN_1135); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1137 = 11'h470 == cnt[10:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1136); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1138 = 11'h471 == cnt[10:0] ? $signed(-32'sh2c27) : $signed(_GEN_1137); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1139 = 11'h472 == cnt[10:0] ? $signed(-32'sh2c8a) : $signed(_GEN_1138); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1140 = 11'h473 == cnt[10:0] ? $signed(-32'sh2ced) : $signed(_GEN_1139); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1141 = 11'h474 == cnt[10:0] ? $signed(-32'sh2d50) : $signed(_GEN_1140); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1142 = 11'h475 == cnt[10:0] ? $signed(-32'sh2db3) : $signed(_GEN_1141); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1143 = 11'h476 == cnt[10:0] ? $signed(-32'sh2e16) : $signed(_GEN_1142); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1144 = 11'h477 == cnt[10:0] ? $signed(-32'sh2e79) : $signed(_GEN_1143); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1145 = 11'h478 == cnt[10:0] ? $signed(-32'sh2edc) : $signed(_GEN_1144); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1146 = 11'h479 == cnt[10:0] ? $signed(-32'sh2f3f) : $signed(_GEN_1145); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1147 = 11'h47a == cnt[10:0] ? $signed(-32'sh2fa1) : $signed(_GEN_1146); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1148 = 11'h47b == cnt[10:0] ? $signed(-32'sh3004) : $signed(_GEN_1147); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1149 = 11'h47c == cnt[10:0] ? $signed(-32'sh3067) : $signed(_GEN_1148); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1150 = 11'h47d == cnt[10:0] ? $signed(-32'sh30ca) : $signed(_GEN_1149); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1151 = 11'h47e == cnt[10:0] ? $signed(-32'sh312c) : $signed(_GEN_1150); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1152 = 11'h47f == cnt[10:0] ? $signed(-32'sh318f) : $signed(_GEN_1151); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1153 = 11'h480 == cnt[10:0] ? $signed(-32'sh31f1) : $signed(_GEN_1152); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1154 = 11'h481 == cnt[10:0] ? $signed(-32'sh3254) : $signed(_GEN_1153); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1155 = 11'h482 == cnt[10:0] ? $signed(-32'sh32b7) : $signed(_GEN_1154); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1156 = 11'h483 == cnt[10:0] ? $signed(-32'sh3319) : $signed(_GEN_1155); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1157 = 11'h484 == cnt[10:0] ? $signed(-32'sh337c) : $signed(_GEN_1156); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1158 = 11'h485 == cnt[10:0] ? $signed(-32'sh33de) : $signed(_GEN_1157); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1159 = 11'h486 == cnt[10:0] ? $signed(-32'sh3440) : $signed(_GEN_1158); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1160 = 11'h487 == cnt[10:0] ? $signed(-32'sh34a3) : $signed(_GEN_1159); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1161 = 11'h488 == cnt[10:0] ? $signed(-32'sh3505) : $signed(_GEN_1160); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1162 = 11'h489 == cnt[10:0] ? $signed(-32'sh3568) : $signed(_GEN_1161); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1163 = 11'h48a == cnt[10:0] ? $signed(-32'sh35ca) : $signed(_GEN_1162); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1164 = 11'h48b == cnt[10:0] ? $signed(-32'sh362c) : $signed(_GEN_1163); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1165 = 11'h48c == cnt[10:0] ? $signed(-32'sh368e) : $signed(_GEN_1164); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1166 = 11'h48d == cnt[10:0] ? $signed(-32'sh36f1) : $signed(_GEN_1165); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1167 = 11'h48e == cnt[10:0] ? $signed(-32'sh3753) : $signed(_GEN_1166); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1168 = 11'h48f == cnt[10:0] ? $signed(-32'sh37b5) : $signed(_GEN_1167); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1169 = 11'h490 == cnt[10:0] ? $signed(-32'sh3817) : $signed(_GEN_1168); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1170 = 11'h491 == cnt[10:0] ? $signed(-32'sh3879) : $signed(_GEN_1169); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1171 = 11'h492 == cnt[10:0] ? $signed(-32'sh38db) : $signed(_GEN_1170); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1172 = 11'h493 == cnt[10:0] ? $signed(-32'sh393d) : $signed(_GEN_1171); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1173 = 11'h494 == cnt[10:0] ? $signed(-32'sh399f) : $signed(_GEN_1172); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1174 = 11'h495 == cnt[10:0] ? $signed(-32'sh3a01) : $signed(_GEN_1173); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1175 = 11'h496 == cnt[10:0] ? $signed(-32'sh3a63) : $signed(_GEN_1174); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1176 = 11'h497 == cnt[10:0] ? $signed(-32'sh3ac5) : $signed(_GEN_1175); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1177 = 11'h498 == cnt[10:0] ? $signed(-32'sh3b27) : $signed(_GEN_1176); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1178 = 11'h499 == cnt[10:0] ? $signed(-32'sh3b88) : $signed(_GEN_1177); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1179 = 11'h49a == cnt[10:0] ? $signed(-32'sh3bea) : $signed(_GEN_1178); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1180 = 11'h49b == cnt[10:0] ? $signed(-32'sh3c4c) : $signed(_GEN_1179); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1181 = 11'h49c == cnt[10:0] ? $signed(-32'sh3cae) : $signed(_GEN_1180); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1182 = 11'h49d == cnt[10:0] ? $signed(-32'sh3d0f) : $signed(_GEN_1181); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1183 = 11'h49e == cnt[10:0] ? $signed(-32'sh3d71) : $signed(_GEN_1182); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1184 = 11'h49f == cnt[10:0] ? $signed(-32'sh3dd2) : $signed(_GEN_1183); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1185 = 11'h4a0 == cnt[10:0] ? $signed(-32'sh3e34) : $signed(_GEN_1184); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1186 = 11'h4a1 == cnt[10:0] ? $signed(-32'sh3e95) : $signed(_GEN_1185); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1187 = 11'h4a2 == cnt[10:0] ? $signed(-32'sh3ef7) : $signed(_GEN_1186); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1188 = 11'h4a3 == cnt[10:0] ? $signed(-32'sh3f58) : $signed(_GEN_1187); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1189 = 11'h4a4 == cnt[10:0] ? $signed(-32'sh3fba) : $signed(_GEN_1188); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1190 = 11'h4a5 == cnt[10:0] ? $signed(-32'sh401b) : $signed(_GEN_1189); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1191 = 11'h4a6 == cnt[10:0] ? $signed(-32'sh407c) : $signed(_GEN_1190); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1192 = 11'h4a7 == cnt[10:0] ? $signed(-32'sh40de) : $signed(_GEN_1191); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1193 = 11'h4a8 == cnt[10:0] ? $signed(-32'sh413f) : $signed(_GEN_1192); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1194 = 11'h4a9 == cnt[10:0] ? $signed(-32'sh41a0) : $signed(_GEN_1193); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1195 = 11'h4aa == cnt[10:0] ? $signed(-32'sh4201) : $signed(_GEN_1194); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1196 = 11'h4ab == cnt[10:0] ? $signed(-32'sh4262) : $signed(_GEN_1195); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1197 = 11'h4ac == cnt[10:0] ? $signed(-32'sh42c3) : $signed(_GEN_1196); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1198 = 11'h4ad == cnt[10:0] ? $signed(-32'sh4324) : $signed(_GEN_1197); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1199 = 11'h4ae == cnt[10:0] ? $signed(-32'sh4385) : $signed(_GEN_1198); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1200 = 11'h4af == cnt[10:0] ? $signed(-32'sh43e6) : $signed(_GEN_1199); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1201 = 11'h4b0 == cnt[10:0] ? $signed(-32'sh4447) : $signed(_GEN_1200); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1202 = 11'h4b1 == cnt[10:0] ? $signed(-32'sh44a8) : $signed(_GEN_1201); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1203 = 11'h4b2 == cnt[10:0] ? $signed(-32'sh4509) : $signed(_GEN_1202); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1204 = 11'h4b3 == cnt[10:0] ? $signed(-32'sh456a) : $signed(_GEN_1203); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1205 = 11'h4b4 == cnt[10:0] ? $signed(-32'sh45cb) : $signed(_GEN_1204); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1206 = 11'h4b5 == cnt[10:0] ? $signed(-32'sh462b) : $signed(_GEN_1205); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1207 = 11'h4b6 == cnt[10:0] ? $signed(-32'sh468c) : $signed(_GEN_1206); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1208 = 11'h4b7 == cnt[10:0] ? $signed(-32'sh46ec) : $signed(_GEN_1207); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1209 = 11'h4b8 == cnt[10:0] ? $signed(-32'sh474d) : $signed(_GEN_1208); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1210 = 11'h4b9 == cnt[10:0] ? $signed(-32'sh47ae) : $signed(_GEN_1209); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1211 = 11'h4ba == cnt[10:0] ? $signed(-32'sh480e) : $signed(_GEN_1210); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1212 = 11'h4bb == cnt[10:0] ? $signed(-32'sh486f) : $signed(_GEN_1211); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1213 = 11'h4bc == cnt[10:0] ? $signed(-32'sh48cf) : $signed(_GEN_1212); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1214 = 11'h4bd == cnt[10:0] ? $signed(-32'sh492f) : $signed(_GEN_1213); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1215 = 11'h4be == cnt[10:0] ? $signed(-32'sh4990) : $signed(_GEN_1214); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1216 = 11'h4bf == cnt[10:0] ? $signed(-32'sh49f0) : $signed(_GEN_1215); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1217 = 11'h4c0 == cnt[10:0] ? $signed(-32'sh4a50) : $signed(_GEN_1216); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1218 = 11'h4c1 == cnt[10:0] ? $signed(-32'sh4ab0) : $signed(_GEN_1217); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1219 = 11'h4c2 == cnt[10:0] ? $signed(-32'sh4b10) : $signed(_GEN_1218); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1220 = 11'h4c3 == cnt[10:0] ? $signed(-32'sh4b71) : $signed(_GEN_1219); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1221 = 11'h4c4 == cnt[10:0] ? $signed(-32'sh4bd1) : $signed(_GEN_1220); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1222 = 11'h4c5 == cnt[10:0] ? $signed(-32'sh4c31) : $signed(_GEN_1221); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1223 = 11'h4c6 == cnt[10:0] ? $signed(-32'sh4c90) : $signed(_GEN_1222); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1224 = 11'h4c7 == cnt[10:0] ? $signed(-32'sh4cf0) : $signed(_GEN_1223); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1225 = 11'h4c8 == cnt[10:0] ? $signed(-32'sh4d50) : $signed(_GEN_1224); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1226 = 11'h4c9 == cnt[10:0] ? $signed(-32'sh4db0) : $signed(_GEN_1225); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1227 = 11'h4ca == cnt[10:0] ? $signed(-32'sh4e10) : $signed(_GEN_1226); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1228 = 11'h4cb == cnt[10:0] ? $signed(-32'sh4e70) : $signed(_GEN_1227); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1229 = 11'h4cc == cnt[10:0] ? $signed(-32'sh4ecf) : $signed(_GEN_1228); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1230 = 11'h4cd == cnt[10:0] ? $signed(-32'sh4f2f) : $signed(_GEN_1229); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1231 = 11'h4ce == cnt[10:0] ? $signed(-32'sh4f8e) : $signed(_GEN_1230); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1232 = 11'h4cf == cnt[10:0] ? $signed(-32'sh4fee) : $signed(_GEN_1231); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1233 = 11'h4d0 == cnt[10:0] ? $signed(-32'sh504d) : $signed(_GEN_1232); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1234 = 11'h4d1 == cnt[10:0] ? $signed(-32'sh50ad) : $signed(_GEN_1233); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1235 = 11'h4d2 == cnt[10:0] ? $signed(-32'sh510c) : $signed(_GEN_1234); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1236 = 11'h4d3 == cnt[10:0] ? $signed(-32'sh516c) : $signed(_GEN_1235); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1237 = 11'h4d4 == cnt[10:0] ? $signed(-32'sh51cb) : $signed(_GEN_1236); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1238 = 11'h4d5 == cnt[10:0] ? $signed(-32'sh522a) : $signed(_GEN_1237); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1239 = 11'h4d6 == cnt[10:0] ? $signed(-32'sh5289) : $signed(_GEN_1238); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1240 = 11'h4d7 == cnt[10:0] ? $signed(-32'sh52e8) : $signed(_GEN_1239); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1241 = 11'h4d8 == cnt[10:0] ? $signed(-32'sh5348) : $signed(_GEN_1240); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1242 = 11'h4d9 == cnt[10:0] ? $signed(-32'sh53a7) : $signed(_GEN_1241); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1243 = 11'h4da == cnt[10:0] ? $signed(-32'sh5406) : $signed(_GEN_1242); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1244 = 11'h4db == cnt[10:0] ? $signed(-32'sh5464) : $signed(_GEN_1243); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1245 = 11'h4dc == cnt[10:0] ? $signed(-32'sh54c3) : $signed(_GEN_1244); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1246 = 11'h4dd == cnt[10:0] ? $signed(-32'sh5522) : $signed(_GEN_1245); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1247 = 11'h4de == cnt[10:0] ? $signed(-32'sh5581) : $signed(_GEN_1246); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1248 = 11'h4df == cnt[10:0] ? $signed(-32'sh55e0) : $signed(_GEN_1247); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1249 = 11'h4e0 == cnt[10:0] ? $signed(-32'sh563e) : $signed(_GEN_1248); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1250 = 11'h4e1 == cnt[10:0] ? $signed(-32'sh569d) : $signed(_GEN_1249); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1251 = 11'h4e2 == cnt[10:0] ? $signed(-32'sh56fc) : $signed(_GEN_1250); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1252 = 11'h4e3 == cnt[10:0] ? $signed(-32'sh575a) : $signed(_GEN_1251); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1253 = 11'h4e4 == cnt[10:0] ? $signed(-32'sh57b9) : $signed(_GEN_1252); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1254 = 11'h4e5 == cnt[10:0] ? $signed(-32'sh5817) : $signed(_GEN_1253); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1255 = 11'h4e6 == cnt[10:0] ? $signed(-32'sh5875) : $signed(_GEN_1254); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1256 = 11'h4e7 == cnt[10:0] ? $signed(-32'sh58d4) : $signed(_GEN_1255); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1257 = 11'h4e8 == cnt[10:0] ? $signed(-32'sh5932) : $signed(_GEN_1256); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1258 = 11'h4e9 == cnt[10:0] ? $signed(-32'sh5990) : $signed(_GEN_1257); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1259 = 11'h4ea == cnt[10:0] ? $signed(-32'sh59ee) : $signed(_GEN_1258); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1260 = 11'h4eb == cnt[10:0] ? $signed(-32'sh5a4c) : $signed(_GEN_1259); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1261 = 11'h4ec == cnt[10:0] ? $signed(-32'sh5aaa) : $signed(_GEN_1260); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1262 = 11'h4ed == cnt[10:0] ? $signed(-32'sh5b08) : $signed(_GEN_1261); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1263 = 11'h4ee == cnt[10:0] ? $signed(-32'sh5b66) : $signed(_GEN_1262); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1264 = 11'h4ef == cnt[10:0] ? $signed(-32'sh5bc4) : $signed(_GEN_1263); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1265 = 11'h4f0 == cnt[10:0] ? $signed(-32'sh5c22) : $signed(_GEN_1264); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1266 = 11'h4f1 == cnt[10:0] ? $signed(-32'sh5c80) : $signed(_GEN_1265); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1267 = 11'h4f2 == cnt[10:0] ? $signed(-32'sh5cde) : $signed(_GEN_1266); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1268 = 11'h4f3 == cnt[10:0] ? $signed(-32'sh5d3b) : $signed(_GEN_1267); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1269 = 11'h4f4 == cnt[10:0] ? $signed(-32'sh5d99) : $signed(_GEN_1268); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1270 = 11'h4f5 == cnt[10:0] ? $signed(-32'sh5df6) : $signed(_GEN_1269); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1271 = 11'h4f6 == cnt[10:0] ? $signed(-32'sh5e54) : $signed(_GEN_1270); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1272 = 11'h4f7 == cnt[10:0] ? $signed(-32'sh5eb1) : $signed(_GEN_1271); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1273 = 11'h4f8 == cnt[10:0] ? $signed(-32'sh5f0f) : $signed(_GEN_1272); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1274 = 11'h4f9 == cnt[10:0] ? $signed(-32'sh5f6c) : $signed(_GEN_1273); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1275 = 11'h4fa == cnt[10:0] ? $signed(-32'sh5fc9) : $signed(_GEN_1274); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1276 = 11'h4fb == cnt[10:0] ? $signed(-32'sh6026) : $signed(_GEN_1275); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1277 = 11'h4fc == cnt[10:0] ? $signed(-32'sh6084) : $signed(_GEN_1276); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1278 = 11'h4fd == cnt[10:0] ? $signed(-32'sh60e1) : $signed(_GEN_1277); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1279 = 11'h4fe == cnt[10:0] ? $signed(-32'sh613e) : $signed(_GEN_1278); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1280 = 11'h4ff == cnt[10:0] ? $signed(-32'sh619b) : $signed(_GEN_1279); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1281 = 11'h500 == cnt[10:0] ? $signed(-32'sh61f8) : $signed(_GEN_1280); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1282 = 11'h501 == cnt[10:0] ? $signed(-32'sh6254) : $signed(_GEN_1281); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1283 = 11'h502 == cnt[10:0] ? $signed(-32'sh62b1) : $signed(_GEN_1282); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1284 = 11'h503 == cnt[10:0] ? $signed(-32'sh630e) : $signed(_GEN_1283); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1285 = 11'h504 == cnt[10:0] ? $signed(-32'sh636b) : $signed(_GEN_1284); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1286 = 11'h505 == cnt[10:0] ? $signed(-32'sh63c7) : $signed(_GEN_1285); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1287 = 11'h506 == cnt[10:0] ? $signed(-32'sh6424) : $signed(_GEN_1286); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1288 = 11'h507 == cnt[10:0] ? $signed(-32'sh6480) : $signed(_GEN_1287); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1289 = 11'h508 == cnt[10:0] ? $signed(-32'sh64dd) : $signed(_GEN_1288); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1290 = 11'h509 == cnt[10:0] ? $signed(-32'sh6539) : $signed(_GEN_1289); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1291 = 11'h50a == cnt[10:0] ? $signed(-32'sh6595) : $signed(_GEN_1290); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1292 = 11'h50b == cnt[10:0] ? $signed(-32'sh65f2) : $signed(_GEN_1291); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1293 = 11'h50c == cnt[10:0] ? $signed(-32'sh664e) : $signed(_GEN_1292); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1294 = 11'h50d == cnt[10:0] ? $signed(-32'sh66aa) : $signed(_GEN_1293); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1295 = 11'h50e == cnt[10:0] ? $signed(-32'sh6706) : $signed(_GEN_1294); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1296 = 11'h50f == cnt[10:0] ? $signed(-32'sh6762) : $signed(_GEN_1295); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1297 = 11'h510 == cnt[10:0] ? $signed(-32'sh67be) : $signed(_GEN_1296); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1298 = 11'h511 == cnt[10:0] ? $signed(-32'sh681a) : $signed(_GEN_1297); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1299 = 11'h512 == cnt[10:0] ? $signed(-32'sh6876) : $signed(_GEN_1298); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1300 = 11'h513 == cnt[10:0] ? $signed(-32'sh68d1) : $signed(_GEN_1299); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1301 = 11'h514 == cnt[10:0] ? $signed(-32'sh692d) : $signed(_GEN_1300); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1302 = 11'h515 == cnt[10:0] ? $signed(-32'sh6989) : $signed(_GEN_1301); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1303 = 11'h516 == cnt[10:0] ? $signed(-32'sh69e4) : $signed(_GEN_1302); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1304 = 11'h517 == cnt[10:0] ? $signed(-32'sh6a40) : $signed(_GEN_1303); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1305 = 11'h518 == cnt[10:0] ? $signed(-32'sh6a9b) : $signed(_GEN_1304); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1306 = 11'h519 == cnt[10:0] ? $signed(-32'sh6af6) : $signed(_GEN_1305); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1307 = 11'h51a == cnt[10:0] ? $signed(-32'sh6b52) : $signed(_GEN_1306); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1308 = 11'h51b == cnt[10:0] ? $signed(-32'sh6bad) : $signed(_GEN_1307); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1309 = 11'h51c == cnt[10:0] ? $signed(-32'sh6c08) : $signed(_GEN_1308); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1310 = 11'h51d == cnt[10:0] ? $signed(-32'sh6c63) : $signed(_GEN_1309); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1311 = 11'h51e == cnt[10:0] ? $signed(-32'sh6cbe) : $signed(_GEN_1310); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1312 = 11'h51f == cnt[10:0] ? $signed(-32'sh6d19) : $signed(_GEN_1311); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1313 = 11'h520 == cnt[10:0] ? $signed(-32'sh6d74) : $signed(_GEN_1312); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1314 = 11'h521 == cnt[10:0] ? $signed(-32'sh6dcf) : $signed(_GEN_1313); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1315 = 11'h522 == cnt[10:0] ? $signed(-32'sh6e2a) : $signed(_GEN_1314); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1316 = 11'h523 == cnt[10:0] ? $signed(-32'sh6e85) : $signed(_GEN_1315); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1317 = 11'h524 == cnt[10:0] ? $signed(-32'sh6edf) : $signed(_GEN_1316); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1318 = 11'h525 == cnt[10:0] ? $signed(-32'sh6f3a) : $signed(_GEN_1317); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1319 = 11'h526 == cnt[10:0] ? $signed(-32'sh6f94) : $signed(_GEN_1318); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1320 = 11'h527 == cnt[10:0] ? $signed(-32'sh6fef) : $signed(_GEN_1319); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1321 = 11'h528 == cnt[10:0] ? $signed(-32'sh7049) : $signed(_GEN_1320); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1322 = 11'h529 == cnt[10:0] ? $signed(-32'sh70a3) : $signed(_GEN_1321); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1323 = 11'h52a == cnt[10:0] ? $signed(-32'sh70fe) : $signed(_GEN_1322); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1324 = 11'h52b == cnt[10:0] ? $signed(-32'sh7158) : $signed(_GEN_1323); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1325 = 11'h52c == cnt[10:0] ? $signed(-32'sh71b2) : $signed(_GEN_1324); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1326 = 11'h52d == cnt[10:0] ? $signed(-32'sh720c) : $signed(_GEN_1325); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1327 = 11'h52e == cnt[10:0] ? $signed(-32'sh7266) : $signed(_GEN_1326); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1328 = 11'h52f == cnt[10:0] ? $signed(-32'sh72c0) : $signed(_GEN_1327); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1329 = 11'h530 == cnt[10:0] ? $signed(-32'sh731a) : $signed(_GEN_1328); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1330 = 11'h531 == cnt[10:0] ? $signed(-32'sh7373) : $signed(_GEN_1329); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1331 = 11'h532 == cnt[10:0] ? $signed(-32'sh73cd) : $signed(_GEN_1330); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1332 = 11'h533 == cnt[10:0] ? $signed(-32'sh7427) : $signed(_GEN_1331); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1333 = 11'h534 == cnt[10:0] ? $signed(-32'sh7480) : $signed(_GEN_1332); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1334 = 11'h535 == cnt[10:0] ? $signed(-32'sh74da) : $signed(_GEN_1333); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1335 = 11'h536 == cnt[10:0] ? $signed(-32'sh7533) : $signed(_GEN_1334); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1336 = 11'h537 == cnt[10:0] ? $signed(-32'sh758d) : $signed(_GEN_1335); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1337 = 11'h538 == cnt[10:0] ? $signed(-32'sh75e6) : $signed(_GEN_1336); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1338 = 11'h539 == cnt[10:0] ? $signed(-32'sh763f) : $signed(_GEN_1337); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1339 = 11'h53a == cnt[10:0] ? $signed(-32'sh7698) : $signed(_GEN_1338); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1340 = 11'h53b == cnt[10:0] ? $signed(-32'sh76f1) : $signed(_GEN_1339); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1341 = 11'h53c == cnt[10:0] ? $signed(-32'sh774a) : $signed(_GEN_1340); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1342 = 11'h53d == cnt[10:0] ? $signed(-32'sh77a3) : $signed(_GEN_1341); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1343 = 11'h53e == cnt[10:0] ? $signed(-32'sh77fc) : $signed(_GEN_1342); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1344 = 11'h53f == cnt[10:0] ? $signed(-32'sh7855) : $signed(_GEN_1343); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1345 = 11'h540 == cnt[10:0] ? $signed(-32'sh78ad) : $signed(_GEN_1344); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1346 = 11'h541 == cnt[10:0] ? $signed(-32'sh7906) : $signed(_GEN_1345); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1347 = 11'h542 == cnt[10:0] ? $signed(-32'sh795f) : $signed(_GEN_1346); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1348 = 11'h543 == cnt[10:0] ? $signed(-32'sh79b7) : $signed(_GEN_1347); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1349 = 11'h544 == cnt[10:0] ? $signed(-32'sh7a10) : $signed(_GEN_1348); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1350 = 11'h545 == cnt[10:0] ? $signed(-32'sh7a68) : $signed(_GEN_1349); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1351 = 11'h546 == cnt[10:0] ? $signed(-32'sh7ac0) : $signed(_GEN_1350); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1352 = 11'h547 == cnt[10:0] ? $signed(-32'sh7b18) : $signed(_GEN_1351); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1353 = 11'h548 == cnt[10:0] ? $signed(-32'sh7b70) : $signed(_GEN_1352); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1354 = 11'h549 == cnt[10:0] ? $signed(-32'sh7bc8) : $signed(_GEN_1353); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1355 = 11'h54a == cnt[10:0] ? $signed(-32'sh7c20) : $signed(_GEN_1354); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1356 = 11'h54b == cnt[10:0] ? $signed(-32'sh7c78) : $signed(_GEN_1355); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1357 = 11'h54c == cnt[10:0] ? $signed(-32'sh7cd0) : $signed(_GEN_1356); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1358 = 11'h54d == cnt[10:0] ? $signed(-32'sh7d28) : $signed(_GEN_1357); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1359 = 11'h54e == cnt[10:0] ? $signed(-32'sh7d7f) : $signed(_GEN_1358); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1360 = 11'h54f == cnt[10:0] ? $signed(-32'sh7dd7) : $signed(_GEN_1359); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1361 = 11'h550 == cnt[10:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1360); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1362 = 11'h551 == cnt[10:0] ? $signed(-32'sh7e86) : $signed(_GEN_1361); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1363 = 11'h552 == cnt[10:0] ? $signed(-32'sh7edd) : $signed(_GEN_1362); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1364 = 11'h553 == cnt[10:0] ? $signed(-32'sh7f35) : $signed(_GEN_1363); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1365 = 11'h554 == cnt[10:0] ? $signed(-32'sh7f8c) : $signed(_GEN_1364); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1366 = 11'h555 == cnt[10:0] ? $signed(-32'sh7fe3) : $signed(_GEN_1365); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1367 = 11'h556 == cnt[10:0] ? $signed(-32'sh803a) : $signed(_GEN_1366); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1368 = 11'h557 == cnt[10:0] ? $signed(-32'sh8091) : $signed(_GEN_1367); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1369 = 11'h558 == cnt[10:0] ? $signed(-32'sh80e8) : $signed(_GEN_1368); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1370 = 11'h559 == cnt[10:0] ? $signed(-32'sh813f) : $signed(_GEN_1369); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1371 = 11'h55a == cnt[10:0] ? $signed(-32'sh8195) : $signed(_GEN_1370); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1372 = 11'h55b == cnt[10:0] ? $signed(-32'sh81ec) : $signed(_GEN_1371); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1373 = 11'h55c == cnt[10:0] ? $signed(-32'sh8243) : $signed(_GEN_1372); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1374 = 11'h55d == cnt[10:0] ? $signed(-32'sh8299) : $signed(_GEN_1373); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1375 = 11'h55e == cnt[10:0] ? $signed(-32'sh82f0) : $signed(_GEN_1374); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1376 = 11'h55f == cnt[10:0] ? $signed(-32'sh8346) : $signed(_GEN_1375); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1377 = 11'h560 == cnt[10:0] ? $signed(-32'sh839c) : $signed(_GEN_1376); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1378 = 11'h561 == cnt[10:0] ? $signed(-32'sh83f2) : $signed(_GEN_1377); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1379 = 11'h562 == cnt[10:0] ? $signed(-32'sh8449) : $signed(_GEN_1378); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1380 = 11'h563 == cnt[10:0] ? $signed(-32'sh849f) : $signed(_GEN_1379); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1381 = 11'h564 == cnt[10:0] ? $signed(-32'sh84f5) : $signed(_GEN_1380); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1382 = 11'h565 == cnt[10:0] ? $signed(-32'sh854a) : $signed(_GEN_1381); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1383 = 11'h566 == cnt[10:0] ? $signed(-32'sh85a0) : $signed(_GEN_1382); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1384 = 11'h567 == cnt[10:0] ? $signed(-32'sh85f6) : $signed(_GEN_1383); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1385 = 11'h568 == cnt[10:0] ? $signed(-32'sh864c) : $signed(_GEN_1384); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1386 = 11'h569 == cnt[10:0] ? $signed(-32'sh86a1) : $signed(_GEN_1385); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1387 = 11'h56a == cnt[10:0] ? $signed(-32'sh86f7) : $signed(_GEN_1386); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1388 = 11'h56b == cnt[10:0] ? $signed(-32'sh874c) : $signed(_GEN_1387); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1389 = 11'h56c == cnt[10:0] ? $signed(-32'sh87a1) : $signed(_GEN_1388); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1390 = 11'h56d == cnt[10:0] ? $signed(-32'sh87f6) : $signed(_GEN_1389); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1391 = 11'h56e == cnt[10:0] ? $signed(-32'sh884c) : $signed(_GEN_1390); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1392 = 11'h56f == cnt[10:0] ? $signed(-32'sh88a1) : $signed(_GEN_1391); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1393 = 11'h570 == cnt[10:0] ? $signed(-32'sh88f6) : $signed(_GEN_1392); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1394 = 11'h571 == cnt[10:0] ? $signed(-32'sh894a) : $signed(_GEN_1393); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1395 = 11'h572 == cnt[10:0] ? $signed(-32'sh899f) : $signed(_GEN_1394); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1396 = 11'h573 == cnt[10:0] ? $signed(-32'sh89f4) : $signed(_GEN_1395); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1397 = 11'h574 == cnt[10:0] ? $signed(-32'sh8a49) : $signed(_GEN_1396); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1398 = 11'h575 == cnt[10:0] ? $signed(-32'sh8a9d) : $signed(_GEN_1397); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1399 = 11'h576 == cnt[10:0] ? $signed(-32'sh8af2) : $signed(_GEN_1398); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1400 = 11'h577 == cnt[10:0] ? $signed(-32'sh8b46) : $signed(_GEN_1399); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1401 = 11'h578 == cnt[10:0] ? $signed(-32'sh8b9a) : $signed(_GEN_1400); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1402 = 11'h579 == cnt[10:0] ? $signed(-32'sh8bef) : $signed(_GEN_1401); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1403 = 11'h57a == cnt[10:0] ? $signed(-32'sh8c43) : $signed(_GEN_1402); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1404 = 11'h57b == cnt[10:0] ? $signed(-32'sh8c97) : $signed(_GEN_1403); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1405 = 11'h57c == cnt[10:0] ? $signed(-32'sh8ceb) : $signed(_GEN_1404); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1406 = 11'h57d == cnt[10:0] ? $signed(-32'sh8d3f) : $signed(_GEN_1405); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1407 = 11'h57e == cnt[10:0] ? $signed(-32'sh8d93) : $signed(_GEN_1406); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1408 = 11'h57f == cnt[10:0] ? $signed(-32'sh8de6) : $signed(_GEN_1407); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1409 = 11'h580 == cnt[10:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1408); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1410 = 11'h581 == cnt[10:0] ? $signed(-32'sh8e8d) : $signed(_GEN_1409); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1411 = 11'h582 == cnt[10:0] ? $signed(-32'sh8ee1) : $signed(_GEN_1410); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1412 = 11'h583 == cnt[10:0] ? $signed(-32'sh8f34) : $signed(_GEN_1411); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1413 = 11'h584 == cnt[10:0] ? $signed(-32'sh8f88) : $signed(_GEN_1412); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1414 = 11'h585 == cnt[10:0] ? $signed(-32'sh8fdb) : $signed(_GEN_1413); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1415 = 11'h586 == cnt[10:0] ? $signed(-32'sh902e) : $signed(_GEN_1414); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1416 = 11'h587 == cnt[10:0] ? $signed(-32'sh9081) : $signed(_GEN_1415); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1417 = 11'h588 == cnt[10:0] ? $signed(-32'sh90d4) : $signed(_GEN_1416); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1418 = 11'h589 == cnt[10:0] ? $signed(-32'sh9127) : $signed(_GEN_1417); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1419 = 11'h58a == cnt[10:0] ? $signed(-32'sh9179) : $signed(_GEN_1418); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1420 = 11'h58b == cnt[10:0] ? $signed(-32'sh91cc) : $signed(_GEN_1419); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1421 = 11'h58c == cnt[10:0] ? $signed(-32'sh921f) : $signed(_GEN_1420); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1422 = 11'h58d == cnt[10:0] ? $signed(-32'sh9271) : $signed(_GEN_1421); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1423 = 11'h58e == cnt[10:0] ? $signed(-32'sh92c4) : $signed(_GEN_1422); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1424 = 11'h58f == cnt[10:0] ? $signed(-32'sh9316) : $signed(_GEN_1423); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1425 = 11'h590 == cnt[10:0] ? $signed(-32'sh9368) : $signed(_GEN_1424); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1426 = 11'h591 == cnt[10:0] ? $signed(-32'sh93ba) : $signed(_GEN_1425); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1427 = 11'h592 == cnt[10:0] ? $signed(-32'sh940c) : $signed(_GEN_1426); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1428 = 11'h593 == cnt[10:0] ? $signed(-32'sh945e) : $signed(_GEN_1427); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1429 = 11'h594 == cnt[10:0] ? $signed(-32'sh94b0) : $signed(_GEN_1428); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1430 = 11'h595 == cnt[10:0] ? $signed(-32'sh9502) : $signed(_GEN_1429); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1431 = 11'h596 == cnt[10:0] ? $signed(-32'sh9554) : $signed(_GEN_1430); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1432 = 11'h597 == cnt[10:0] ? $signed(-32'sh95a5) : $signed(_GEN_1431); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1433 = 11'h598 == cnt[10:0] ? $signed(-32'sh95f7) : $signed(_GEN_1432); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1434 = 11'h599 == cnt[10:0] ? $signed(-32'sh9648) : $signed(_GEN_1433); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1435 = 11'h59a == cnt[10:0] ? $signed(-32'sh969a) : $signed(_GEN_1434); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1436 = 11'h59b == cnt[10:0] ? $signed(-32'sh96eb) : $signed(_GEN_1435); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1437 = 11'h59c == cnt[10:0] ? $signed(-32'sh973c) : $signed(_GEN_1436); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1438 = 11'h59d == cnt[10:0] ? $signed(-32'sh978d) : $signed(_GEN_1437); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1439 = 11'h59e == cnt[10:0] ? $signed(-32'sh97de) : $signed(_GEN_1438); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1440 = 11'h59f == cnt[10:0] ? $signed(-32'sh982f) : $signed(_GEN_1439); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1441 = 11'h5a0 == cnt[10:0] ? $signed(-32'sh9880) : $signed(_GEN_1440); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1442 = 11'h5a1 == cnt[10:0] ? $signed(-32'sh98d0) : $signed(_GEN_1441); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1443 = 11'h5a2 == cnt[10:0] ? $signed(-32'sh9921) : $signed(_GEN_1442); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1444 = 11'h5a3 == cnt[10:0] ? $signed(-32'sh9972) : $signed(_GEN_1443); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1445 = 11'h5a4 == cnt[10:0] ? $signed(-32'sh99c2) : $signed(_GEN_1444); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1446 = 11'h5a5 == cnt[10:0] ? $signed(-32'sh9a12) : $signed(_GEN_1445); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1447 = 11'h5a6 == cnt[10:0] ? $signed(-32'sh9a63) : $signed(_GEN_1446); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1448 = 11'h5a7 == cnt[10:0] ? $signed(-32'sh9ab3) : $signed(_GEN_1447); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1449 = 11'h5a8 == cnt[10:0] ? $signed(-32'sh9b03) : $signed(_GEN_1448); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1450 = 11'h5a9 == cnt[10:0] ? $signed(-32'sh9b53) : $signed(_GEN_1449); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1451 = 11'h5aa == cnt[10:0] ? $signed(-32'sh9ba3) : $signed(_GEN_1450); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1452 = 11'h5ab == cnt[10:0] ? $signed(-32'sh9bf2) : $signed(_GEN_1451); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1453 = 11'h5ac == cnt[10:0] ? $signed(-32'sh9c42) : $signed(_GEN_1452); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1454 = 11'h5ad == cnt[10:0] ? $signed(-32'sh9c92) : $signed(_GEN_1453); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1455 = 11'h5ae == cnt[10:0] ? $signed(-32'sh9ce1) : $signed(_GEN_1454); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1456 = 11'h5af == cnt[10:0] ? $signed(-32'sh9d31) : $signed(_GEN_1455); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1457 = 11'h5b0 == cnt[10:0] ? $signed(-32'sh9d80) : $signed(_GEN_1456); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1458 = 11'h5b1 == cnt[10:0] ? $signed(-32'sh9dcf) : $signed(_GEN_1457); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1459 = 11'h5b2 == cnt[10:0] ? $signed(-32'sh9e1e) : $signed(_GEN_1458); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1460 = 11'h5b3 == cnt[10:0] ? $signed(-32'sh9e6d) : $signed(_GEN_1459); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1461 = 11'h5b4 == cnt[10:0] ? $signed(-32'sh9ebc) : $signed(_GEN_1460); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1462 = 11'h5b5 == cnt[10:0] ? $signed(-32'sh9f0b) : $signed(_GEN_1461); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1463 = 11'h5b6 == cnt[10:0] ? $signed(-32'sh9f5a) : $signed(_GEN_1462); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1464 = 11'h5b7 == cnt[10:0] ? $signed(-32'sh9fa8) : $signed(_GEN_1463); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1465 = 11'h5b8 == cnt[10:0] ? $signed(-32'sh9ff7) : $signed(_GEN_1464); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1466 = 11'h5b9 == cnt[10:0] ? $signed(-32'sha045) : $signed(_GEN_1465); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1467 = 11'h5ba == cnt[10:0] ? $signed(-32'sha094) : $signed(_GEN_1466); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1468 = 11'h5bb == cnt[10:0] ? $signed(-32'sha0e2) : $signed(_GEN_1467); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1469 = 11'h5bc == cnt[10:0] ? $signed(-32'sha130) : $signed(_GEN_1468); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1470 = 11'h5bd == cnt[10:0] ? $signed(-32'sha17e) : $signed(_GEN_1469); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1471 = 11'h5be == cnt[10:0] ? $signed(-32'sha1cc) : $signed(_GEN_1470); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1472 = 11'h5bf == cnt[10:0] ? $signed(-32'sha21a) : $signed(_GEN_1471); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1473 = 11'h5c0 == cnt[10:0] ? $signed(-32'sha268) : $signed(_GEN_1472); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1474 = 11'h5c1 == cnt[10:0] ? $signed(-32'sha2b5) : $signed(_GEN_1473); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1475 = 11'h5c2 == cnt[10:0] ? $signed(-32'sha303) : $signed(_GEN_1474); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1476 = 11'h5c3 == cnt[10:0] ? $signed(-32'sha350) : $signed(_GEN_1475); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1477 = 11'h5c4 == cnt[10:0] ? $signed(-32'sha39e) : $signed(_GEN_1476); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1478 = 11'h5c5 == cnt[10:0] ? $signed(-32'sha3eb) : $signed(_GEN_1477); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1479 = 11'h5c6 == cnt[10:0] ? $signed(-32'sha438) : $signed(_GEN_1478); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1480 = 11'h5c7 == cnt[10:0] ? $signed(-32'sha485) : $signed(_GEN_1479); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1481 = 11'h5c8 == cnt[10:0] ? $signed(-32'sha4d2) : $signed(_GEN_1480); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1482 = 11'h5c9 == cnt[10:0] ? $signed(-32'sha51f) : $signed(_GEN_1481); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1483 = 11'h5ca == cnt[10:0] ? $signed(-32'sha56c) : $signed(_GEN_1482); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1484 = 11'h5cb == cnt[10:0] ? $signed(-32'sha5b8) : $signed(_GEN_1483); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1485 = 11'h5cc == cnt[10:0] ? $signed(-32'sha605) : $signed(_GEN_1484); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1486 = 11'h5cd == cnt[10:0] ? $signed(-32'sha652) : $signed(_GEN_1485); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1487 = 11'h5ce == cnt[10:0] ? $signed(-32'sha69e) : $signed(_GEN_1486); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1488 = 11'h5cf == cnt[10:0] ? $signed(-32'sha6ea) : $signed(_GEN_1487); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1489 = 11'h5d0 == cnt[10:0] ? $signed(-32'sha736) : $signed(_GEN_1488); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1490 = 11'h5d1 == cnt[10:0] ? $signed(-32'sha782) : $signed(_GEN_1489); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1491 = 11'h5d2 == cnt[10:0] ? $signed(-32'sha7ce) : $signed(_GEN_1490); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1492 = 11'h5d3 == cnt[10:0] ? $signed(-32'sha81a) : $signed(_GEN_1491); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1493 = 11'h5d4 == cnt[10:0] ? $signed(-32'sha866) : $signed(_GEN_1492); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1494 = 11'h5d5 == cnt[10:0] ? $signed(-32'sha8b2) : $signed(_GEN_1493); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1495 = 11'h5d6 == cnt[10:0] ? $signed(-32'sha8fd) : $signed(_GEN_1494); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1496 = 11'h5d7 == cnt[10:0] ? $signed(-32'sha949) : $signed(_GEN_1495); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1497 = 11'h5d8 == cnt[10:0] ? $signed(-32'sha994) : $signed(_GEN_1496); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1498 = 11'h5d9 == cnt[10:0] ? $signed(-32'sha9df) : $signed(_GEN_1497); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1499 = 11'h5da == cnt[10:0] ? $signed(-32'shaa2a) : $signed(_GEN_1498); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1500 = 11'h5db == cnt[10:0] ? $signed(-32'shaa76) : $signed(_GEN_1499); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1501 = 11'h5dc == cnt[10:0] ? $signed(-32'shaac1) : $signed(_GEN_1500); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1502 = 11'h5dd == cnt[10:0] ? $signed(-32'shab0b) : $signed(_GEN_1501); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1503 = 11'h5de == cnt[10:0] ? $signed(-32'shab56) : $signed(_GEN_1502); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1504 = 11'h5df == cnt[10:0] ? $signed(-32'shaba1) : $signed(_GEN_1503); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1505 = 11'h5e0 == cnt[10:0] ? $signed(-32'shabeb) : $signed(_GEN_1504); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1506 = 11'h5e1 == cnt[10:0] ? $signed(-32'shac36) : $signed(_GEN_1505); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1507 = 11'h5e2 == cnt[10:0] ? $signed(-32'shac80) : $signed(_GEN_1506); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1508 = 11'h5e3 == cnt[10:0] ? $signed(-32'shacca) : $signed(_GEN_1507); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1509 = 11'h5e4 == cnt[10:0] ? $signed(-32'shad14) : $signed(_GEN_1508); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1510 = 11'h5e5 == cnt[10:0] ? $signed(-32'shad5e) : $signed(_GEN_1509); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1511 = 11'h5e6 == cnt[10:0] ? $signed(-32'shada8) : $signed(_GEN_1510); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1512 = 11'h5e7 == cnt[10:0] ? $signed(-32'shadf2) : $signed(_GEN_1511); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1513 = 11'h5e8 == cnt[10:0] ? $signed(-32'shae3c) : $signed(_GEN_1512); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1514 = 11'h5e9 == cnt[10:0] ? $signed(-32'shae85) : $signed(_GEN_1513); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1515 = 11'h5ea == cnt[10:0] ? $signed(-32'shaecf) : $signed(_GEN_1514); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1516 = 11'h5eb == cnt[10:0] ? $signed(-32'shaf18) : $signed(_GEN_1515); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1517 = 11'h5ec == cnt[10:0] ? $signed(-32'shaf62) : $signed(_GEN_1516); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1518 = 11'h5ed == cnt[10:0] ? $signed(-32'shafab) : $signed(_GEN_1517); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1519 = 11'h5ee == cnt[10:0] ? $signed(-32'shaff4) : $signed(_GEN_1518); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1520 = 11'h5ef == cnt[10:0] ? $signed(-32'shb03d) : $signed(_GEN_1519); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1521 = 11'h5f0 == cnt[10:0] ? $signed(-32'shb086) : $signed(_GEN_1520); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1522 = 11'h5f1 == cnt[10:0] ? $signed(-32'shb0ce) : $signed(_GEN_1521); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1523 = 11'h5f2 == cnt[10:0] ? $signed(-32'shb117) : $signed(_GEN_1522); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1524 = 11'h5f3 == cnt[10:0] ? $signed(-32'shb160) : $signed(_GEN_1523); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1525 = 11'h5f4 == cnt[10:0] ? $signed(-32'shb1a8) : $signed(_GEN_1524); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1526 = 11'h5f5 == cnt[10:0] ? $signed(-32'shb1f0) : $signed(_GEN_1525); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1527 = 11'h5f6 == cnt[10:0] ? $signed(-32'shb239) : $signed(_GEN_1526); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1528 = 11'h5f7 == cnt[10:0] ? $signed(-32'shb281) : $signed(_GEN_1527); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1529 = 11'h5f8 == cnt[10:0] ? $signed(-32'shb2c9) : $signed(_GEN_1528); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1530 = 11'h5f9 == cnt[10:0] ? $signed(-32'shb311) : $signed(_GEN_1529); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1531 = 11'h5fa == cnt[10:0] ? $signed(-32'shb358) : $signed(_GEN_1530); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1532 = 11'h5fb == cnt[10:0] ? $signed(-32'shb3a0) : $signed(_GEN_1531); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1533 = 11'h5fc == cnt[10:0] ? $signed(-32'shb3e8) : $signed(_GEN_1532); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1534 = 11'h5fd == cnt[10:0] ? $signed(-32'shb42f) : $signed(_GEN_1533); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1535 = 11'h5fe == cnt[10:0] ? $signed(-32'shb477) : $signed(_GEN_1534); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1536 = 11'h5ff == cnt[10:0] ? $signed(-32'shb4be) : $signed(_GEN_1535); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1537 = 11'h600 == cnt[10:0] ? $signed(-32'shb505) : $signed(_GEN_1536); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1538 = 11'h601 == cnt[10:0] ? $signed(-32'shb54c) : $signed(_GEN_1537); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1539 = 11'h602 == cnt[10:0] ? $signed(-32'shb593) : $signed(_GEN_1538); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1540 = 11'h603 == cnt[10:0] ? $signed(-32'shb5da) : $signed(_GEN_1539); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1541 = 11'h604 == cnt[10:0] ? $signed(-32'shb620) : $signed(_GEN_1540); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1542 = 11'h605 == cnt[10:0] ? $signed(-32'shb667) : $signed(_GEN_1541); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1543 = 11'h606 == cnt[10:0] ? $signed(-32'shb6ad) : $signed(_GEN_1542); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1544 = 11'h607 == cnt[10:0] ? $signed(-32'shb6f4) : $signed(_GEN_1543); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1545 = 11'h608 == cnt[10:0] ? $signed(-32'shb73a) : $signed(_GEN_1544); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1546 = 11'h609 == cnt[10:0] ? $signed(-32'shb780) : $signed(_GEN_1545); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1547 = 11'h60a == cnt[10:0] ? $signed(-32'shb7c6) : $signed(_GEN_1546); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1548 = 11'h60b == cnt[10:0] ? $signed(-32'shb80c) : $signed(_GEN_1547); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1549 = 11'h60c == cnt[10:0] ? $signed(-32'shb852) : $signed(_GEN_1548); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1550 = 11'h60d == cnt[10:0] ? $signed(-32'shb898) : $signed(_GEN_1549); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1551 = 11'h60e == cnt[10:0] ? $signed(-32'shb8dd) : $signed(_GEN_1550); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1552 = 11'h60f == cnt[10:0] ? $signed(-32'shb923) : $signed(_GEN_1551); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1553 = 11'h610 == cnt[10:0] ? $signed(-32'shb968) : $signed(_GEN_1552); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1554 = 11'h611 == cnt[10:0] ? $signed(-32'shb9ae) : $signed(_GEN_1553); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1555 = 11'h612 == cnt[10:0] ? $signed(-32'shb9f3) : $signed(_GEN_1554); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1556 = 11'h613 == cnt[10:0] ? $signed(-32'shba38) : $signed(_GEN_1555); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1557 = 11'h614 == cnt[10:0] ? $signed(-32'shba7d) : $signed(_GEN_1556); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1558 = 11'h615 == cnt[10:0] ? $signed(-32'shbac1) : $signed(_GEN_1557); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1559 = 11'h616 == cnt[10:0] ? $signed(-32'shbb06) : $signed(_GEN_1558); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1560 = 11'h617 == cnt[10:0] ? $signed(-32'shbb4b) : $signed(_GEN_1559); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1561 = 11'h618 == cnt[10:0] ? $signed(-32'shbb8f) : $signed(_GEN_1560); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1562 = 11'h619 == cnt[10:0] ? $signed(-32'shbbd4) : $signed(_GEN_1561); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1563 = 11'h61a == cnt[10:0] ? $signed(-32'shbc18) : $signed(_GEN_1562); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1564 = 11'h61b == cnt[10:0] ? $signed(-32'shbc5c) : $signed(_GEN_1563); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1565 = 11'h61c == cnt[10:0] ? $signed(-32'shbca0) : $signed(_GEN_1564); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1566 = 11'h61d == cnt[10:0] ? $signed(-32'shbce4) : $signed(_GEN_1565); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1567 = 11'h61e == cnt[10:0] ? $signed(-32'shbd28) : $signed(_GEN_1566); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1568 = 11'h61f == cnt[10:0] ? $signed(-32'shbd6b) : $signed(_GEN_1567); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1569 = 11'h620 == cnt[10:0] ? $signed(-32'shbdaf) : $signed(_GEN_1568); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1570 = 11'h621 == cnt[10:0] ? $signed(-32'shbdf2) : $signed(_GEN_1569); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1571 = 11'h622 == cnt[10:0] ? $signed(-32'shbe36) : $signed(_GEN_1570); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1572 = 11'h623 == cnt[10:0] ? $signed(-32'shbe79) : $signed(_GEN_1571); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1573 = 11'h624 == cnt[10:0] ? $signed(-32'shbebc) : $signed(_GEN_1572); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1574 = 11'h625 == cnt[10:0] ? $signed(-32'shbeff) : $signed(_GEN_1573); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1575 = 11'h626 == cnt[10:0] ? $signed(-32'shbf42) : $signed(_GEN_1574); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1576 = 11'h627 == cnt[10:0] ? $signed(-32'shbf85) : $signed(_GEN_1575); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1577 = 11'h628 == cnt[10:0] ? $signed(-32'shbfc7) : $signed(_GEN_1576); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1578 = 11'h629 == cnt[10:0] ? $signed(-32'shc00a) : $signed(_GEN_1577); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1579 = 11'h62a == cnt[10:0] ? $signed(-32'shc04c) : $signed(_GEN_1578); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1580 = 11'h62b == cnt[10:0] ? $signed(-32'shc08f) : $signed(_GEN_1579); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1581 = 11'h62c == cnt[10:0] ? $signed(-32'shc0d1) : $signed(_GEN_1580); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1582 = 11'h62d == cnt[10:0] ? $signed(-32'shc113) : $signed(_GEN_1581); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1583 = 11'h62e == cnt[10:0] ? $signed(-32'shc155) : $signed(_GEN_1582); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1584 = 11'h62f == cnt[10:0] ? $signed(-32'shc197) : $signed(_GEN_1583); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1585 = 11'h630 == cnt[10:0] ? $signed(-32'shc1d8) : $signed(_GEN_1584); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1586 = 11'h631 == cnt[10:0] ? $signed(-32'shc21a) : $signed(_GEN_1585); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1587 = 11'h632 == cnt[10:0] ? $signed(-32'shc25c) : $signed(_GEN_1586); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1588 = 11'h633 == cnt[10:0] ? $signed(-32'shc29d) : $signed(_GEN_1587); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1589 = 11'h634 == cnt[10:0] ? $signed(-32'shc2de) : $signed(_GEN_1588); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1590 = 11'h635 == cnt[10:0] ? $signed(-32'shc31f) : $signed(_GEN_1589); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1591 = 11'h636 == cnt[10:0] ? $signed(-32'shc360) : $signed(_GEN_1590); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1592 = 11'h637 == cnt[10:0] ? $signed(-32'shc3a1) : $signed(_GEN_1591); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1593 = 11'h638 == cnt[10:0] ? $signed(-32'shc3e2) : $signed(_GEN_1592); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1594 = 11'h639 == cnt[10:0] ? $signed(-32'shc423) : $signed(_GEN_1593); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1595 = 11'h63a == cnt[10:0] ? $signed(-32'shc463) : $signed(_GEN_1594); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1596 = 11'h63b == cnt[10:0] ? $signed(-32'shc4a4) : $signed(_GEN_1595); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1597 = 11'h63c == cnt[10:0] ? $signed(-32'shc4e4) : $signed(_GEN_1596); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1598 = 11'h63d == cnt[10:0] ? $signed(-32'shc524) : $signed(_GEN_1597); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1599 = 11'h63e == cnt[10:0] ? $signed(-32'shc564) : $signed(_GEN_1598); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1600 = 11'h63f == cnt[10:0] ? $signed(-32'shc5a4) : $signed(_GEN_1599); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1601 = 11'h640 == cnt[10:0] ? $signed(-32'shc5e4) : $signed(_GEN_1600); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1602 = 11'h641 == cnt[10:0] ? $signed(-32'shc624) : $signed(_GEN_1601); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1603 = 11'h642 == cnt[10:0] ? $signed(-32'shc663) : $signed(_GEN_1602); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1604 = 11'h643 == cnt[10:0] ? $signed(-32'shc6a3) : $signed(_GEN_1603); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1605 = 11'h644 == cnt[10:0] ? $signed(-32'shc6e2) : $signed(_GEN_1604); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1606 = 11'h645 == cnt[10:0] ? $signed(-32'shc721) : $signed(_GEN_1605); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1607 = 11'h646 == cnt[10:0] ? $signed(-32'shc761) : $signed(_GEN_1606); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1608 = 11'h647 == cnt[10:0] ? $signed(-32'shc7a0) : $signed(_GEN_1607); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1609 = 11'h648 == cnt[10:0] ? $signed(-32'shc7de) : $signed(_GEN_1608); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1610 = 11'h649 == cnt[10:0] ? $signed(-32'shc81d) : $signed(_GEN_1609); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1611 = 11'h64a == cnt[10:0] ? $signed(-32'shc85c) : $signed(_GEN_1610); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1612 = 11'h64b == cnt[10:0] ? $signed(-32'shc89a) : $signed(_GEN_1611); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1613 = 11'h64c == cnt[10:0] ? $signed(-32'shc8d9) : $signed(_GEN_1612); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1614 = 11'h64d == cnt[10:0] ? $signed(-32'shc917) : $signed(_GEN_1613); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1615 = 11'h64e == cnt[10:0] ? $signed(-32'shc955) : $signed(_GEN_1614); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1616 = 11'h64f == cnt[10:0] ? $signed(-32'shc993) : $signed(_GEN_1615); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1617 = 11'h650 == cnt[10:0] ? $signed(-32'shc9d1) : $signed(_GEN_1616); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1618 = 11'h651 == cnt[10:0] ? $signed(-32'shca0f) : $signed(_GEN_1617); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1619 = 11'h652 == cnt[10:0] ? $signed(-32'shca4d) : $signed(_GEN_1618); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1620 = 11'h653 == cnt[10:0] ? $signed(-32'shca8a) : $signed(_GEN_1619); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1621 = 11'h654 == cnt[10:0] ? $signed(-32'shcac7) : $signed(_GEN_1620); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1622 = 11'h655 == cnt[10:0] ? $signed(-32'shcb05) : $signed(_GEN_1621); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1623 = 11'h656 == cnt[10:0] ? $signed(-32'shcb42) : $signed(_GEN_1622); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1624 = 11'h657 == cnt[10:0] ? $signed(-32'shcb7f) : $signed(_GEN_1623); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1625 = 11'h658 == cnt[10:0] ? $signed(-32'shcbbc) : $signed(_GEN_1624); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1626 = 11'h659 == cnt[10:0] ? $signed(-32'shcbf9) : $signed(_GEN_1625); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1627 = 11'h65a == cnt[10:0] ? $signed(-32'shcc35) : $signed(_GEN_1626); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1628 = 11'h65b == cnt[10:0] ? $signed(-32'shcc72) : $signed(_GEN_1627); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1629 = 11'h65c == cnt[10:0] ? $signed(-32'shccae) : $signed(_GEN_1628); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1630 = 11'h65d == cnt[10:0] ? $signed(-32'shcceb) : $signed(_GEN_1629); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1631 = 11'h65e == cnt[10:0] ? $signed(-32'shcd27) : $signed(_GEN_1630); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1632 = 11'h65f == cnt[10:0] ? $signed(-32'shcd63) : $signed(_GEN_1631); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1633 = 11'h660 == cnt[10:0] ? $signed(-32'shcd9f) : $signed(_GEN_1632); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1634 = 11'h661 == cnt[10:0] ? $signed(-32'shcddb) : $signed(_GEN_1633); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1635 = 11'h662 == cnt[10:0] ? $signed(-32'shce17) : $signed(_GEN_1634); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1636 = 11'h663 == cnt[10:0] ? $signed(-32'shce52) : $signed(_GEN_1635); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1637 = 11'h664 == cnt[10:0] ? $signed(-32'shce8e) : $signed(_GEN_1636); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1638 = 11'h665 == cnt[10:0] ? $signed(-32'shcec9) : $signed(_GEN_1637); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1639 = 11'h666 == cnt[10:0] ? $signed(-32'shcf04) : $signed(_GEN_1638); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1640 = 11'h667 == cnt[10:0] ? $signed(-32'shcf3f) : $signed(_GEN_1639); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1641 = 11'h668 == cnt[10:0] ? $signed(-32'shcf7a) : $signed(_GEN_1640); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1642 = 11'h669 == cnt[10:0] ? $signed(-32'shcfb5) : $signed(_GEN_1641); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1643 = 11'h66a == cnt[10:0] ? $signed(-32'shcff0) : $signed(_GEN_1642); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1644 = 11'h66b == cnt[10:0] ? $signed(-32'shd02a) : $signed(_GEN_1643); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1645 = 11'h66c == cnt[10:0] ? $signed(-32'shd065) : $signed(_GEN_1644); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1646 = 11'h66d == cnt[10:0] ? $signed(-32'shd09f) : $signed(_GEN_1645); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1647 = 11'h66e == cnt[10:0] ? $signed(-32'shd0d9) : $signed(_GEN_1646); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1648 = 11'h66f == cnt[10:0] ? $signed(-32'shd113) : $signed(_GEN_1647); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1649 = 11'h670 == cnt[10:0] ? $signed(-32'shd14d) : $signed(_GEN_1648); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1650 = 11'h671 == cnt[10:0] ? $signed(-32'shd187) : $signed(_GEN_1649); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1651 = 11'h672 == cnt[10:0] ? $signed(-32'shd1c1) : $signed(_GEN_1650); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1652 = 11'h673 == cnt[10:0] ? $signed(-32'shd1fa) : $signed(_GEN_1651); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1653 = 11'h674 == cnt[10:0] ? $signed(-32'shd234) : $signed(_GEN_1652); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1654 = 11'h675 == cnt[10:0] ? $signed(-32'shd26d) : $signed(_GEN_1653); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1655 = 11'h676 == cnt[10:0] ? $signed(-32'shd2a6) : $signed(_GEN_1654); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1656 = 11'h677 == cnt[10:0] ? $signed(-32'shd2df) : $signed(_GEN_1655); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1657 = 11'h678 == cnt[10:0] ? $signed(-32'shd318) : $signed(_GEN_1656); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1658 = 11'h679 == cnt[10:0] ? $signed(-32'shd351) : $signed(_GEN_1657); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1659 = 11'h67a == cnt[10:0] ? $signed(-32'shd38a) : $signed(_GEN_1658); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1660 = 11'h67b == cnt[10:0] ? $signed(-32'shd3c2) : $signed(_GEN_1659); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1661 = 11'h67c == cnt[10:0] ? $signed(-32'shd3fb) : $signed(_GEN_1660); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1662 = 11'h67d == cnt[10:0] ? $signed(-32'shd433) : $signed(_GEN_1661); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1663 = 11'h67e == cnt[10:0] ? $signed(-32'shd46b) : $signed(_GEN_1662); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1664 = 11'h67f == cnt[10:0] ? $signed(-32'shd4a3) : $signed(_GEN_1663); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1665 = 11'h680 == cnt[10:0] ? $signed(-32'shd4db) : $signed(_GEN_1664); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1666 = 11'h681 == cnt[10:0] ? $signed(-32'shd513) : $signed(_GEN_1665); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1667 = 11'h682 == cnt[10:0] ? $signed(-32'shd54b) : $signed(_GEN_1666); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1668 = 11'h683 == cnt[10:0] ? $signed(-32'shd582) : $signed(_GEN_1667); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1669 = 11'h684 == cnt[10:0] ? $signed(-32'shd5ba) : $signed(_GEN_1668); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1670 = 11'h685 == cnt[10:0] ? $signed(-32'shd5f1) : $signed(_GEN_1669); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1671 = 11'h686 == cnt[10:0] ? $signed(-32'shd628) : $signed(_GEN_1670); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1672 = 11'h687 == cnt[10:0] ? $signed(-32'shd65f) : $signed(_GEN_1671); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1673 = 11'h688 == cnt[10:0] ? $signed(-32'shd696) : $signed(_GEN_1672); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1674 = 11'h689 == cnt[10:0] ? $signed(-32'shd6cd) : $signed(_GEN_1673); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1675 = 11'h68a == cnt[10:0] ? $signed(-32'shd703) : $signed(_GEN_1674); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1676 = 11'h68b == cnt[10:0] ? $signed(-32'shd73a) : $signed(_GEN_1675); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1677 = 11'h68c == cnt[10:0] ? $signed(-32'shd770) : $signed(_GEN_1676); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1678 = 11'h68d == cnt[10:0] ? $signed(-32'shd7a6) : $signed(_GEN_1677); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1679 = 11'h68e == cnt[10:0] ? $signed(-32'shd7dc) : $signed(_GEN_1678); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1680 = 11'h68f == cnt[10:0] ? $signed(-32'shd812) : $signed(_GEN_1679); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1681 = 11'h690 == cnt[10:0] ? $signed(-32'shd848) : $signed(_GEN_1680); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1682 = 11'h691 == cnt[10:0] ? $signed(-32'shd87e) : $signed(_GEN_1681); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1683 = 11'h692 == cnt[10:0] ? $signed(-32'shd8b4) : $signed(_GEN_1682); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1684 = 11'h693 == cnt[10:0] ? $signed(-32'shd8e9) : $signed(_GEN_1683); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1685 = 11'h694 == cnt[10:0] ? $signed(-32'shd91e) : $signed(_GEN_1684); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1686 = 11'h695 == cnt[10:0] ? $signed(-32'shd954) : $signed(_GEN_1685); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1687 = 11'h696 == cnt[10:0] ? $signed(-32'shd989) : $signed(_GEN_1686); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1688 = 11'h697 == cnt[10:0] ? $signed(-32'shd9be) : $signed(_GEN_1687); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1689 = 11'h698 == cnt[10:0] ? $signed(-32'shd9f2) : $signed(_GEN_1688); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1690 = 11'h699 == cnt[10:0] ? $signed(-32'shda27) : $signed(_GEN_1689); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1691 = 11'h69a == cnt[10:0] ? $signed(-32'shda5c) : $signed(_GEN_1690); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1692 = 11'h69b == cnt[10:0] ? $signed(-32'shda90) : $signed(_GEN_1691); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1693 = 11'h69c == cnt[10:0] ? $signed(-32'shdac4) : $signed(_GEN_1692); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1694 = 11'h69d == cnt[10:0] ? $signed(-32'shdaf8) : $signed(_GEN_1693); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1695 = 11'h69e == cnt[10:0] ? $signed(-32'shdb2c) : $signed(_GEN_1694); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1696 = 11'h69f == cnt[10:0] ? $signed(-32'shdb60) : $signed(_GEN_1695); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1697 = 11'h6a0 == cnt[10:0] ? $signed(-32'shdb94) : $signed(_GEN_1696); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1698 = 11'h6a1 == cnt[10:0] ? $signed(-32'shdbc8) : $signed(_GEN_1697); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1699 = 11'h6a2 == cnt[10:0] ? $signed(-32'shdbfb) : $signed(_GEN_1698); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1700 = 11'h6a3 == cnt[10:0] ? $signed(-32'shdc2f) : $signed(_GEN_1699); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1701 = 11'h6a4 == cnt[10:0] ? $signed(-32'shdc62) : $signed(_GEN_1700); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1702 = 11'h6a5 == cnt[10:0] ? $signed(-32'shdc95) : $signed(_GEN_1701); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1703 = 11'h6a6 == cnt[10:0] ? $signed(-32'shdcc8) : $signed(_GEN_1702); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1704 = 11'h6a7 == cnt[10:0] ? $signed(-32'shdcfb) : $signed(_GEN_1703); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1705 = 11'h6a8 == cnt[10:0] ? $signed(-32'shdd2d) : $signed(_GEN_1704); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1706 = 11'h6a9 == cnt[10:0] ? $signed(-32'shdd60) : $signed(_GEN_1705); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1707 = 11'h6aa == cnt[10:0] ? $signed(-32'shdd92) : $signed(_GEN_1706); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1708 = 11'h6ab == cnt[10:0] ? $signed(-32'shddc5) : $signed(_GEN_1707); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1709 = 11'h6ac == cnt[10:0] ? $signed(-32'shddf7) : $signed(_GEN_1708); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1710 = 11'h6ad == cnt[10:0] ? $signed(-32'shde29) : $signed(_GEN_1709); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1711 = 11'h6ae == cnt[10:0] ? $signed(-32'shde5b) : $signed(_GEN_1710); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1712 = 11'h6af == cnt[10:0] ? $signed(-32'shde8c) : $signed(_GEN_1711); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1713 = 11'h6b0 == cnt[10:0] ? $signed(-32'shdebe) : $signed(_GEN_1712); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1714 = 11'h6b1 == cnt[10:0] ? $signed(-32'shdef0) : $signed(_GEN_1713); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1715 = 11'h6b2 == cnt[10:0] ? $signed(-32'shdf21) : $signed(_GEN_1714); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1716 = 11'h6b3 == cnt[10:0] ? $signed(-32'shdf52) : $signed(_GEN_1715); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1717 = 11'h6b4 == cnt[10:0] ? $signed(-32'shdf83) : $signed(_GEN_1716); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1718 = 11'h6b5 == cnt[10:0] ? $signed(-32'shdfb4) : $signed(_GEN_1717); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1719 = 11'h6b6 == cnt[10:0] ? $signed(-32'shdfe5) : $signed(_GEN_1718); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1720 = 11'h6b7 == cnt[10:0] ? $signed(-32'she016) : $signed(_GEN_1719); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1721 = 11'h6b8 == cnt[10:0] ? $signed(-32'she046) : $signed(_GEN_1720); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1722 = 11'h6b9 == cnt[10:0] ? $signed(-32'she077) : $signed(_GEN_1721); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1723 = 11'h6ba == cnt[10:0] ? $signed(-32'she0a7) : $signed(_GEN_1722); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1724 = 11'h6bb == cnt[10:0] ? $signed(-32'she0d7) : $signed(_GEN_1723); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1725 = 11'h6bc == cnt[10:0] ? $signed(-32'she107) : $signed(_GEN_1724); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1726 = 11'h6bd == cnt[10:0] ? $signed(-32'she137) : $signed(_GEN_1725); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1727 = 11'h6be == cnt[10:0] ? $signed(-32'she167) : $signed(_GEN_1726); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1728 = 11'h6bf == cnt[10:0] ? $signed(-32'she196) : $signed(_GEN_1727); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1729 = 11'h6c0 == cnt[10:0] ? $signed(-32'she1c6) : $signed(_GEN_1728); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1730 = 11'h6c1 == cnt[10:0] ? $signed(-32'she1f5) : $signed(_GEN_1729); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1731 = 11'h6c2 == cnt[10:0] ? $signed(-32'she224) : $signed(_GEN_1730); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1732 = 11'h6c3 == cnt[10:0] ? $signed(-32'she253) : $signed(_GEN_1731); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1733 = 11'h6c4 == cnt[10:0] ? $signed(-32'she282) : $signed(_GEN_1732); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1734 = 11'h6c5 == cnt[10:0] ? $signed(-32'she2b1) : $signed(_GEN_1733); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1735 = 11'h6c6 == cnt[10:0] ? $signed(-32'she2df) : $signed(_GEN_1734); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1736 = 11'h6c7 == cnt[10:0] ? $signed(-32'she30e) : $signed(_GEN_1735); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1737 = 11'h6c8 == cnt[10:0] ? $signed(-32'she33c) : $signed(_GEN_1736); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1738 = 11'h6c9 == cnt[10:0] ? $signed(-32'she36b) : $signed(_GEN_1737); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1739 = 11'h6ca == cnt[10:0] ? $signed(-32'she399) : $signed(_GEN_1738); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1740 = 11'h6cb == cnt[10:0] ? $signed(-32'she3c7) : $signed(_GEN_1739); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1741 = 11'h6cc == cnt[10:0] ? $signed(-32'she3f4) : $signed(_GEN_1740); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1742 = 11'h6cd == cnt[10:0] ? $signed(-32'she422) : $signed(_GEN_1741); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1743 = 11'h6ce == cnt[10:0] ? $signed(-32'she450) : $signed(_GEN_1742); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1744 = 11'h6cf == cnt[10:0] ? $signed(-32'she47d) : $signed(_GEN_1743); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1745 = 11'h6d0 == cnt[10:0] ? $signed(-32'she4aa) : $signed(_GEN_1744); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1746 = 11'h6d1 == cnt[10:0] ? $signed(-32'she4d7) : $signed(_GEN_1745); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1747 = 11'h6d2 == cnt[10:0] ? $signed(-32'she504) : $signed(_GEN_1746); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1748 = 11'h6d3 == cnt[10:0] ? $signed(-32'she531) : $signed(_GEN_1747); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1749 = 11'h6d4 == cnt[10:0] ? $signed(-32'she55e) : $signed(_GEN_1748); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1750 = 11'h6d5 == cnt[10:0] ? $signed(-32'she58b) : $signed(_GEN_1749); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1751 = 11'h6d6 == cnt[10:0] ? $signed(-32'she5b7) : $signed(_GEN_1750); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1752 = 11'h6d7 == cnt[10:0] ? $signed(-32'she5e3) : $signed(_GEN_1751); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1753 = 11'h6d8 == cnt[10:0] ? $signed(-32'she610) : $signed(_GEN_1752); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1754 = 11'h6d9 == cnt[10:0] ? $signed(-32'she63c) : $signed(_GEN_1753); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1755 = 11'h6da == cnt[10:0] ? $signed(-32'she667) : $signed(_GEN_1754); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1756 = 11'h6db == cnt[10:0] ? $signed(-32'she693) : $signed(_GEN_1755); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1757 = 11'h6dc == cnt[10:0] ? $signed(-32'she6bf) : $signed(_GEN_1756); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1758 = 11'h6dd == cnt[10:0] ? $signed(-32'she6ea) : $signed(_GEN_1757); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1759 = 11'h6de == cnt[10:0] ? $signed(-32'she716) : $signed(_GEN_1758); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1760 = 11'h6df == cnt[10:0] ? $signed(-32'she741) : $signed(_GEN_1759); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1761 = 11'h6e0 == cnt[10:0] ? $signed(-32'she76c) : $signed(_GEN_1760); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1762 = 11'h6e1 == cnt[10:0] ? $signed(-32'she797) : $signed(_GEN_1761); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1763 = 11'h6e2 == cnt[10:0] ? $signed(-32'she7c2) : $signed(_GEN_1762); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1764 = 11'h6e3 == cnt[10:0] ? $signed(-32'she7ec) : $signed(_GEN_1763); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1765 = 11'h6e4 == cnt[10:0] ? $signed(-32'she817) : $signed(_GEN_1764); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1766 = 11'h6e5 == cnt[10:0] ? $signed(-32'she841) : $signed(_GEN_1765); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1767 = 11'h6e6 == cnt[10:0] ? $signed(-32'she86b) : $signed(_GEN_1766); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1768 = 11'h6e7 == cnt[10:0] ? $signed(-32'she895) : $signed(_GEN_1767); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1769 = 11'h6e8 == cnt[10:0] ? $signed(-32'she8bf) : $signed(_GEN_1768); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1770 = 11'h6e9 == cnt[10:0] ? $signed(-32'she8e9) : $signed(_GEN_1769); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1771 = 11'h6ea == cnt[10:0] ? $signed(-32'she913) : $signed(_GEN_1770); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1772 = 11'h6eb == cnt[10:0] ? $signed(-32'she93c) : $signed(_GEN_1771); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1773 = 11'h6ec == cnt[10:0] ? $signed(-32'she966) : $signed(_GEN_1772); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1774 = 11'h6ed == cnt[10:0] ? $signed(-32'she98f) : $signed(_GEN_1773); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1775 = 11'h6ee == cnt[10:0] ? $signed(-32'she9b8) : $signed(_GEN_1774); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1776 = 11'h6ef == cnt[10:0] ? $signed(-32'she9e1) : $signed(_GEN_1775); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1777 = 11'h6f0 == cnt[10:0] ? $signed(-32'shea0a) : $signed(_GEN_1776); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1778 = 11'h6f1 == cnt[10:0] ? $signed(-32'shea32) : $signed(_GEN_1777); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1779 = 11'h6f2 == cnt[10:0] ? $signed(-32'shea5b) : $signed(_GEN_1778); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1780 = 11'h6f3 == cnt[10:0] ? $signed(-32'shea83) : $signed(_GEN_1779); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1781 = 11'h6f4 == cnt[10:0] ? $signed(-32'sheaab) : $signed(_GEN_1780); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1782 = 11'h6f5 == cnt[10:0] ? $signed(-32'shead4) : $signed(_GEN_1781); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1783 = 11'h6f6 == cnt[10:0] ? $signed(-32'sheafc) : $signed(_GEN_1782); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1784 = 11'h6f7 == cnt[10:0] ? $signed(-32'sheb23) : $signed(_GEN_1783); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1785 = 11'h6f8 == cnt[10:0] ? $signed(-32'sheb4b) : $signed(_GEN_1784); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1786 = 11'h6f9 == cnt[10:0] ? $signed(-32'sheb73) : $signed(_GEN_1785); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1787 = 11'h6fa == cnt[10:0] ? $signed(-32'sheb9a) : $signed(_GEN_1786); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1788 = 11'h6fb == cnt[10:0] ? $signed(-32'shebc1) : $signed(_GEN_1787); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1789 = 11'h6fc == cnt[10:0] ? $signed(-32'shebe8) : $signed(_GEN_1788); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1790 = 11'h6fd == cnt[10:0] ? $signed(-32'shec0f) : $signed(_GEN_1789); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1791 = 11'h6fe == cnt[10:0] ? $signed(-32'shec36) : $signed(_GEN_1790); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1792 = 11'h6ff == cnt[10:0] ? $signed(-32'shec5d) : $signed(_GEN_1791); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1793 = 11'h700 == cnt[10:0] ? $signed(-32'shec83) : $signed(_GEN_1792); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1794 = 11'h701 == cnt[10:0] ? $signed(-32'shecaa) : $signed(_GEN_1793); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1795 = 11'h702 == cnt[10:0] ? $signed(-32'shecd0) : $signed(_GEN_1794); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1796 = 11'h703 == cnt[10:0] ? $signed(-32'shecf6) : $signed(_GEN_1795); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1797 = 11'h704 == cnt[10:0] ? $signed(-32'shed1c) : $signed(_GEN_1796); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1798 = 11'h705 == cnt[10:0] ? $signed(-32'shed42) : $signed(_GEN_1797); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1799 = 11'h706 == cnt[10:0] ? $signed(-32'shed68) : $signed(_GEN_1798); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1800 = 11'h707 == cnt[10:0] ? $signed(-32'shed8d) : $signed(_GEN_1799); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1801 = 11'h708 == cnt[10:0] ? $signed(-32'shedb3) : $signed(_GEN_1800); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1802 = 11'h709 == cnt[10:0] ? $signed(-32'shedd8) : $signed(_GEN_1801); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1803 = 11'h70a == cnt[10:0] ? $signed(-32'shedfd) : $signed(_GEN_1802); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1804 = 11'h70b == cnt[10:0] ? $signed(-32'shee22) : $signed(_GEN_1803); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1805 = 11'h70c == cnt[10:0] ? $signed(-32'shee47) : $signed(_GEN_1804); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1806 = 11'h70d == cnt[10:0] ? $signed(-32'shee6b) : $signed(_GEN_1805); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1807 = 11'h70e == cnt[10:0] ? $signed(-32'shee90) : $signed(_GEN_1806); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1808 = 11'h70f == cnt[10:0] ? $signed(-32'sheeb4) : $signed(_GEN_1807); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1809 = 11'h710 == cnt[10:0] ? $signed(-32'sheed9) : $signed(_GEN_1808); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1810 = 11'h711 == cnt[10:0] ? $signed(-32'sheefd) : $signed(_GEN_1809); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1811 = 11'h712 == cnt[10:0] ? $signed(-32'shef21) : $signed(_GEN_1810); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1812 = 11'h713 == cnt[10:0] ? $signed(-32'shef45) : $signed(_GEN_1811); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1813 = 11'h714 == cnt[10:0] ? $signed(-32'shef68) : $signed(_GEN_1812); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1814 = 11'h715 == cnt[10:0] ? $signed(-32'shef8c) : $signed(_GEN_1813); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1815 = 11'h716 == cnt[10:0] ? $signed(-32'shefaf) : $signed(_GEN_1814); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1816 = 11'h717 == cnt[10:0] ? $signed(-32'shefd2) : $signed(_GEN_1815); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1817 = 11'h718 == cnt[10:0] ? $signed(-32'sheff5) : $signed(_GEN_1816); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1818 = 11'h719 == cnt[10:0] ? $signed(-32'shf018) : $signed(_GEN_1817); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1819 = 11'h71a == cnt[10:0] ? $signed(-32'shf03b) : $signed(_GEN_1818); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1820 = 11'h71b == cnt[10:0] ? $signed(-32'shf05e) : $signed(_GEN_1819); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1821 = 11'h71c == cnt[10:0] ? $signed(-32'shf080) : $signed(_GEN_1820); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1822 = 11'h71d == cnt[10:0] ? $signed(-32'shf0a3) : $signed(_GEN_1821); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1823 = 11'h71e == cnt[10:0] ? $signed(-32'shf0c5) : $signed(_GEN_1822); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1824 = 11'h71f == cnt[10:0] ? $signed(-32'shf0e7) : $signed(_GEN_1823); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1825 = 11'h720 == cnt[10:0] ? $signed(-32'shf109) : $signed(_GEN_1824); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1826 = 11'h721 == cnt[10:0] ? $signed(-32'shf12b) : $signed(_GEN_1825); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1827 = 11'h722 == cnt[10:0] ? $signed(-32'shf14c) : $signed(_GEN_1826); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1828 = 11'h723 == cnt[10:0] ? $signed(-32'shf16e) : $signed(_GEN_1827); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1829 = 11'h724 == cnt[10:0] ? $signed(-32'shf18f) : $signed(_GEN_1828); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1830 = 11'h725 == cnt[10:0] ? $signed(-32'shf1b1) : $signed(_GEN_1829); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1831 = 11'h726 == cnt[10:0] ? $signed(-32'shf1d2) : $signed(_GEN_1830); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1832 = 11'h727 == cnt[10:0] ? $signed(-32'shf1f3) : $signed(_GEN_1831); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1833 = 11'h728 == cnt[10:0] ? $signed(-32'shf213) : $signed(_GEN_1832); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1834 = 11'h729 == cnt[10:0] ? $signed(-32'shf234) : $signed(_GEN_1833); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1835 = 11'h72a == cnt[10:0] ? $signed(-32'shf254) : $signed(_GEN_1834); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1836 = 11'h72b == cnt[10:0] ? $signed(-32'shf275) : $signed(_GEN_1835); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1837 = 11'h72c == cnt[10:0] ? $signed(-32'shf295) : $signed(_GEN_1836); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1838 = 11'h72d == cnt[10:0] ? $signed(-32'shf2b5) : $signed(_GEN_1837); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1839 = 11'h72e == cnt[10:0] ? $signed(-32'shf2d5) : $signed(_GEN_1838); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1840 = 11'h72f == cnt[10:0] ? $signed(-32'shf2f5) : $signed(_GEN_1839); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1841 = 11'h730 == cnt[10:0] ? $signed(-32'shf314) : $signed(_GEN_1840); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1842 = 11'h731 == cnt[10:0] ? $signed(-32'shf334) : $signed(_GEN_1841); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1843 = 11'h732 == cnt[10:0] ? $signed(-32'shf353) : $signed(_GEN_1842); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1844 = 11'h733 == cnt[10:0] ? $signed(-32'shf372) : $signed(_GEN_1843); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1845 = 11'h734 == cnt[10:0] ? $signed(-32'shf391) : $signed(_GEN_1844); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1846 = 11'h735 == cnt[10:0] ? $signed(-32'shf3b0) : $signed(_GEN_1845); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1847 = 11'h736 == cnt[10:0] ? $signed(-32'shf3cf) : $signed(_GEN_1846); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1848 = 11'h737 == cnt[10:0] ? $signed(-32'shf3ed) : $signed(_GEN_1847); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1849 = 11'h738 == cnt[10:0] ? $signed(-32'shf40c) : $signed(_GEN_1848); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1850 = 11'h739 == cnt[10:0] ? $signed(-32'shf42a) : $signed(_GEN_1849); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1851 = 11'h73a == cnt[10:0] ? $signed(-32'shf448) : $signed(_GEN_1850); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1852 = 11'h73b == cnt[10:0] ? $signed(-32'shf466) : $signed(_GEN_1851); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1853 = 11'h73c == cnt[10:0] ? $signed(-32'shf484) : $signed(_GEN_1852); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1854 = 11'h73d == cnt[10:0] ? $signed(-32'shf4a2) : $signed(_GEN_1853); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1855 = 11'h73e == cnt[10:0] ? $signed(-32'shf4bf) : $signed(_GEN_1854); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1856 = 11'h73f == cnt[10:0] ? $signed(-32'shf4dd) : $signed(_GEN_1855); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1857 = 11'h740 == cnt[10:0] ? $signed(-32'shf4fa) : $signed(_GEN_1856); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1858 = 11'h741 == cnt[10:0] ? $signed(-32'shf517) : $signed(_GEN_1857); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1859 = 11'h742 == cnt[10:0] ? $signed(-32'shf534) : $signed(_GEN_1858); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1860 = 11'h743 == cnt[10:0] ? $signed(-32'shf551) : $signed(_GEN_1859); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1861 = 11'h744 == cnt[10:0] ? $signed(-32'shf56e) : $signed(_GEN_1860); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1862 = 11'h745 == cnt[10:0] ? $signed(-32'shf58a) : $signed(_GEN_1861); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1863 = 11'h746 == cnt[10:0] ? $signed(-32'shf5a6) : $signed(_GEN_1862); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1864 = 11'h747 == cnt[10:0] ? $signed(-32'shf5c3) : $signed(_GEN_1863); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1865 = 11'h748 == cnt[10:0] ? $signed(-32'shf5df) : $signed(_GEN_1864); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1866 = 11'h749 == cnt[10:0] ? $signed(-32'shf5fb) : $signed(_GEN_1865); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1867 = 11'h74a == cnt[10:0] ? $signed(-32'shf616) : $signed(_GEN_1866); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1868 = 11'h74b == cnt[10:0] ? $signed(-32'shf632) : $signed(_GEN_1867); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1869 = 11'h74c == cnt[10:0] ? $signed(-32'shf64e) : $signed(_GEN_1868); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1870 = 11'h74d == cnt[10:0] ? $signed(-32'shf669) : $signed(_GEN_1869); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1871 = 11'h74e == cnt[10:0] ? $signed(-32'shf684) : $signed(_GEN_1870); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1872 = 11'h74f == cnt[10:0] ? $signed(-32'shf69f) : $signed(_GEN_1871); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1873 = 11'h750 == cnt[10:0] ? $signed(-32'shf6ba) : $signed(_GEN_1872); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1874 = 11'h751 == cnt[10:0] ? $signed(-32'shf6d5) : $signed(_GEN_1873); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1875 = 11'h752 == cnt[10:0] ? $signed(-32'shf6ef) : $signed(_GEN_1874); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1876 = 11'h753 == cnt[10:0] ? $signed(-32'shf70a) : $signed(_GEN_1875); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1877 = 11'h754 == cnt[10:0] ? $signed(-32'shf724) : $signed(_GEN_1876); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1878 = 11'h755 == cnt[10:0] ? $signed(-32'shf73e) : $signed(_GEN_1877); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1879 = 11'h756 == cnt[10:0] ? $signed(-32'shf758) : $signed(_GEN_1878); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1880 = 11'h757 == cnt[10:0] ? $signed(-32'shf772) : $signed(_GEN_1879); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1881 = 11'h758 == cnt[10:0] ? $signed(-32'shf78c) : $signed(_GEN_1880); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1882 = 11'h759 == cnt[10:0] ? $signed(-32'shf7a5) : $signed(_GEN_1881); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1883 = 11'h75a == cnt[10:0] ? $signed(-32'shf7bf) : $signed(_GEN_1882); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1884 = 11'h75b == cnt[10:0] ? $signed(-32'shf7d8) : $signed(_GEN_1883); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1885 = 11'h75c == cnt[10:0] ? $signed(-32'shf7f1) : $signed(_GEN_1884); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1886 = 11'h75d == cnt[10:0] ? $signed(-32'shf80a) : $signed(_GEN_1885); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1887 = 11'h75e == cnt[10:0] ? $signed(-32'shf823) : $signed(_GEN_1886); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1888 = 11'h75f == cnt[10:0] ? $signed(-32'shf83b) : $signed(_GEN_1887); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1889 = 11'h760 == cnt[10:0] ? $signed(-32'shf854) : $signed(_GEN_1888); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1890 = 11'h761 == cnt[10:0] ? $signed(-32'shf86c) : $signed(_GEN_1889); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1891 = 11'h762 == cnt[10:0] ? $signed(-32'shf885) : $signed(_GEN_1890); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1892 = 11'h763 == cnt[10:0] ? $signed(-32'shf89d) : $signed(_GEN_1891); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1893 = 11'h764 == cnt[10:0] ? $signed(-32'shf8b4) : $signed(_GEN_1892); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1894 = 11'h765 == cnt[10:0] ? $signed(-32'shf8cc) : $signed(_GEN_1893); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1895 = 11'h766 == cnt[10:0] ? $signed(-32'shf8e4) : $signed(_GEN_1894); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1896 = 11'h767 == cnt[10:0] ? $signed(-32'shf8fb) : $signed(_GEN_1895); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1897 = 11'h768 == cnt[10:0] ? $signed(-32'shf913) : $signed(_GEN_1896); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1898 = 11'h769 == cnt[10:0] ? $signed(-32'shf92a) : $signed(_GEN_1897); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1899 = 11'h76a == cnt[10:0] ? $signed(-32'shf941) : $signed(_GEN_1898); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1900 = 11'h76b == cnt[10:0] ? $signed(-32'shf958) : $signed(_GEN_1899); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1901 = 11'h76c == cnt[10:0] ? $signed(-32'shf96e) : $signed(_GEN_1900); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1902 = 11'h76d == cnt[10:0] ? $signed(-32'shf985) : $signed(_GEN_1901); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1903 = 11'h76e == cnt[10:0] ? $signed(-32'shf99b) : $signed(_GEN_1902); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1904 = 11'h76f == cnt[10:0] ? $signed(-32'shf9b2) : $signed(_GEN_1903); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1905 = 11'h770 == cnt[10:0] ? $signed(-32'shf9c8) : $signed(_GEN_1904); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1906 = 11'h771 == cnt[10:0] ? $signed(-32'shf9de) : $signed(_GEN_1905); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1907 = 11'h772 == cnt[10:0] ? $signed(-32'shf9f3) : $signed(_GEN_1906); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1908 = 11'h773 == cnt[10:0] ? $signed(-32'shfa09) : $signed(_GEN_1907); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1909 = 11'h774 == cnt[10:0] ? $signed(-32'shfa1f) : $signed(_GEN_1908); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1910 = 11'h775 == cnt[10:0] ? $signed(-32'shfa34) : $signed(_GEN_1909); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1911 = 11'h776 == cnt[10:0] ? $signed(-32'shfa49) : $signed(_GEN_1910); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1912 = 11'h777 == cnt[10:0] ? $signed(-32'shfa5e) : $signed(_GEN_1911); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1913 = 11'h778 == cnt[10:0] ? $signed(-32'shfa73) : $signed(_GEN_1912); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1914 = 11'h779 == cnt[10:0] ? $signed(-32'shfa88) : $signed(_GEN_1913); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1915 = 11'h77a == cnt[10:0] ? $signed(-32'shfa9c) : $signed(_GEN_1914); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1916 = 11'h77b == cnt[10:0] ? $signed(-32'shfab1) : $signed(_GEN_1915); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1917 = 11'h77c == cnt[10:0] ? $signed(-32'shfac5) : $signed(_GEN_1916); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1918 = 11'h77d == cnt[10:0] ? $signed(-32'shfad9) : $signed(_GEN_1917); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1919 = 11'h77e == cnt[10:0] ? $signed(-32'shfaed) : $signed(_GEN_1918); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1920 = 11'h77f == cnt[10:0] ? $signed(-32'shfb01) : $signed(_GEN_1919); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1921 = 11'h780 == cnt[10:0] ? $signed(-32'shfb15) : $signed(_GEN_1920); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1922 = 11'h781 == cnt[10:0] ? $signed(-32'shfb28) : $signed(_GEN_1921); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1923 = 11'h782 == cnt[10:0] ? $signed(-32'shfb3c) : $signed(_GEN_1922); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1924 = 11'h783 == cnt[10:0] ? $signed(-32'shfb4f) : $signed(_GEN_1923); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1925 = 11'h784 == cnt[10:0] ? $signed(-32'shfb62) : $signed(_GEN_1924); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1926 = 11'h785 == cnt[10:0] ? $signed(-32'shfb75) : $signed(_GEN_1925); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1927 = 11'h786 == cnt[10:0] ? $signed(-32'shfb88) : $signed(_GEN_1926); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1928 = 11'h787 == cnt[10:0] ? $signed(-32'shfb9a) : $signed(_GEN_1927); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1929 = 11'h788 == cnt[10:0] ? $signed(-32'shfbad) : $signed(_GEN_1928); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1930 = 11'h789 == cnt[10:0] ? $signed(-32'shfbbf) : $signed(_GEN_1929); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1931 = 11'h78a == cnt[10:0] ? $signed(-32'shfbd1) : $signed(_GEN_1930); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1932 = 11'h78b == cnt[10:0] ? $signed(-32'shfbe3) : $signed(_GEN_1931); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1933 = 11'h78c == cnt[10:0] ? $signed(-32'shfbf5) : $signed(_GEN_1932); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1934 = 11'h78d == cnt[10:0] ? $signed(-32'shfc07) : $signed(_GEN_1933); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1935 = 11'h78e == cnt[10:0] ? $signed(-32'shfc18) : $signed(_GEN_1934); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1936 = 11'h78f == cnt[10:0] ? $signed(-32'shfc2a) : $signed(_GEN_1935); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1937 = 11'h790 == cnt[10:0] ? $signed(-32'shfc3b) : $signed(_GEN_1936); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1938 = 11'h791 == cnt[10:0] ? $signed(-32'shfc4c) : $signed(_GEN_1937); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1939 = 11'h792 == cnt[10:0] ? $signed(-32'shfc5d) : $signed(_GEN_1938); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1940 = 11'h793 == cnt[10:0] ? $signed(-32'shfc6e) : $signed(_GEN_1939); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1941 = 11'h794 == cnt[10:0] ? $signed(-32'shfc7f) : $signed(_GEN_1940); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1942 = 11'h795 == cnt[10:0] ? $signed(-32'shfc8f) : $signed(_GEN_1941); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1943 = 11'h796 == cnt[10:0] ? $signed(-32'shfca0) : $signed(_GEN_1942); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1944 = 11'h797 == cnt[10:0] ? $signed(-32'shfcb0) : $signed(_GEN_1943); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1945 = 11'h798 == cnt[10:0] ? $signed(-32'shfcc0) : $signed(_GEN_1944); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1946 = 11'h799 == cnt[10:0] ? $signed(-32'shfcd0) : $signed(_GEN_1945); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1947 = 11'h79a == cnt[10:0] ? $signed(-32'shfcdf) : $signed(_GEN_1946); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1948 = 11'h79b == cnt[10:0] ? $signed(-32'shfcef) : $signed(_GEN_1947); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1949 = 11'h79c == cnt[10:0] ? $signed(-32'shfcfe) : $signed(_GEN_1948); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1950 = 11'h79d == cnt[10:0] ? $signed(-32'shfd0e) : $signed(_GEN_1949); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1951 = 11'h79e == cnt[10:0] ? $signed(-32'shfd1d) : $signed(_GEN_1950); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1952 = 11'h79f == cnt[10:0] ? $signed(-32'shfd2c) : $signed(_GEN_1951); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1953 = 11'h7a0 == cnt[10:0] ? $signed(-32'shfd3b) : $signed(_GEN_1952); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1954 = 11'h7a1 == cnt[10:0] ? $signed(-32'shfd49) : $signed(_GEN_1953); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1955 = 11'h7a2 == cnt[10:0] ? $signed(-32'shfd58) : $signed(_GEN_1954); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1956 = 11'h7a3 == cnt[10:0] ? $signed(-32'shfd66) : $signed(_GEN_1955); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1957 = 11'h7a4 == cnt[10:0] ? $signed(-32'shfd74) : $signed(_GEN_1956); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1958 = 11'h7a5 == cnt[10:0] ? $signed(-32'shfd83) : $signed(_GEN_1957); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1959 = 11'h7a6 == cnt[10:0] ? $signed(-32'shfd90) : $signed(_GEN_1958); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1960 = 11'h7a7 == cnt[10:0] ? $signed(-32'shfd9e) : $signed(_GEN_1959); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1961 = 11'h7a8 == cnt[10:0] ? $signed(-32'shfdac) : $signed(_GEN_1960); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1962 = 11'h7a9 == cnt[10:0] ? $signed(-32'shfdb9) : $signed(_GEN_1961); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1963 = 11'h7aa == cnt[10:0] ? $signed(-32'shfdc7) : $signed(_GEN_1962); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1964 = 11'h7ab == cnt[10:0] ? $signed(-32'shfdd4) : $signed(_GEN_1963); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1965 = 11'h7ac == cnt[10:0] ? $signed(-32'shfde1) : $signed(_GEN_1964); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1966 = 11'h7ad == cnt[10:0] ? $signed(-32'shfdee) : $signed(_GEN_1965); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1967 = 11'h7ae == cnt[10:0] ? $signed(-32'shfdfa) : $signed(_GEN_1966); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1968 = 11'h7af == cnt[10:0] ? $signed(-32'shfe07) : $signed(_GEN_1967); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1969 = 11'h7b0 == cnt[10:0] ? $signed(-32'shfe13) : $signed(_GEN_1968); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1970 = 11'h7b1 == cnt[10:0] ? $signed(-32'shfe1f) : $signed(_GEN_1969); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1971 = 11'h7b2 == cnt[10:0] ? $signed(-32'shfe2b) : $signed(_GEN_1970); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1972 = 11'h7b3 == cnt[10:0] ? $signed(-32'shfe37) : $signed(_GEN_1971); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1973 = 11'h7b4 == cnt[10:0] ? $signed(-32'shfe43) : $signed(_GEN_1972); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1974 = 11'h7b5 == cnt[10:0] ? $signed(-32'shfe4f) : $signed(_GEN_1973); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1975 = 11'h7b6 == cnt[10:0] ? $signed(-32'shfe5a) : $signed(_GEN_1974); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1976 = 11'h7b7 == cnt[10:0] ? $signed(-32'shfe66) : $signed(_GEN_1975); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1977 = 11'h7b8 == cnt[10:0] ? $signed(-32'shfe71) : $signed(_GEN_1976); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1978 = 11'h7b9 == cnt[10:0] ? $signed(-32'shfe7c) : $signed(_GEN_1977); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1979 = 11'h7ba == cnt[10:0] ? $signed(-32'shfe87) : $signed(_GEN_1978); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1980 = 11'h7bb == cnt[10:0] ? $signed(-32'shfe91) : $signed(_GEN_1979); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1981 = 11'h7bc == cnt[10:0] ? $signed(-32'shfe9c) : $signed(_GEN_1980); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1982 = 11'h7bd == cnt[10:0] ? $signed(-32'shfea6) : $signed(_GEN_1981); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1983 = 11'h7be == cnt[10:0] ? $signed(-32'shfeb0) : $signed(_GEN_1982); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1984 = 11'h7bf == cnt[10:0] ? $signed(-32'shfeba) : $signed(_GEN_1983); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1985 = 11'h7c0 == cnt[10:0] ? $signed(-32'shfec4) : $signed(_GEN_1984); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1986 = 11'h7c1 == cnt[10:0] ? $signed(-32'shfece) : $signed(_GEN_1985); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1987 = 11'h7c2 == cnt[10:0] ? $signed(-32'shfed8) : $signed(_GEN_1986); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1988 = 11'h7c3 == cnt[10:0] ? $signed(-32'shfee1) : $signed(_GEN_1987); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1989 = 11'h7c4 == cnt[10:0] ? $signed(-32'shfeeb) : $signed(_GEN_1988); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1990 = 11'h7c5 == cnt[10:0] ? $signed(-32'shfef4) : $signed(_GEN_1989); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1991 = 11'h7c6 == cnt[10:0] ? $signed(-32'shfefd) : $signed(_GEN_1990); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1992 = 11'h7c7 == cnt[10:0] ? $signed(-32'shff06) : $signed(_GEN_1991); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1993 = 11'h7c8 == cnt[10:0] ? $signed(-32'shff0e) : $signed(_GEN_1992); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1994 = 11'h7c9 == cnt[10:0] ? $signed(-32'shff17) : $signed(_GEN_1993); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1995 = 11'h7ca == cnt[10:0] ? $signed(-32'shff1f) : $signed(_GEN_1994); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1996 = 11'h7cb == cnt[10:0] ? $signed(-32'shff28) : $signed(_GEN_1995); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1997 = 11'h7cc == cnt[10:0] ? $signed(-32'shff30) : $signed(_GEN_1996); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1998 = 11'h7cd == cnt[10:0] ? $signed(-32'shff38) : $signed(_GEN_1997); // @[FFT.scala 34:12]
  wire [31:0] _GEN_1999 = 11'h7ce == cnt[10:0] ? $signed(-32'shff3f) : $signed(_GEN_1998); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2000 = 11'h7cf == cnt[10:0] ? $signed(-32'shff47) : $signed(_GEN_1999); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2001 = 11'h7d0 == cnt[10:0] ? $signed(-32'shff4e) : $signed(_GEN_2000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2002 = 11'h7d1 == cnt[10:0] ? $signed(-32'shff56) : $signed(_GEN_2001); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2003 = 11'h7d2 == cnt[10:0] ? $signed(-32'shff5d) : $signed(_GEN_2002); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2004 = 11'h7d3 == cnt[10:0] ? $signed(-32'shff64) : $signed(_GEN_2003); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2005 = 11'h7d4 == cnt[10:0] ? $signed(-32'shff6b) : $signed(_GEN_2004); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2006 = 11'h7d5 == cnt[10:0] ? $signed(-32'shff71) : $signed(_GEN_2005); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2007 = 11'h7d6 == cnt[10:0] ? $signed(-32'shff78) : $signed(_GEN_2006); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2008 = 11'h7d7 == cnt[10:0] ? $signed(-32'shff7e) : $signed(_GEN_2007); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2009 = 11'h7d8 == cnt[10:0] ? $signed(-32'shff85) : $signed(_GEN_2008); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2010 = 11'h7d9 == cnt[10:0] ? $signed(-32'shff8b) : $signed(_GEN_2009); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2011 = 11'h7da == cnt[10:0] ? $signed(-32'shff91) : $signed(_GEN_2010); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2012 = 11'h7db == cnt[10:0] ? $signed(-32'shff96) : $signed(_GEN_2011); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2013 = 11'h7dc == cnt[10:0] ? $signed(-32'shff9c) : $signed(_GEN_2012); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2014 = 11'h7dd == cnt[10:0] ? $signed(-32'shffa2) : $signed(_GEN_2013); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2015 = 11'h7de == cnt[10:0] ? $signed(-32'shffa7) : $signed(_GEN_2014); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2016 = 11'h7df == cnt[10:0] ? $signed(-32'shffac) : $signed(_GEN_2015); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2017 = 11'h7e0 == cnt[10:0] ? $signed(-32'shffb1) : $signed(_GEN_2016); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2018 = 11'h7e1 == cnt[10:0] ? $signed(-32'shffb6) : $signed(_GEN_2017); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2019 = 11'h7e2 == cnt[10:0] ? $signed(-32'shffbb) : $signed(_GEN_2018); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2020 = 11'h7e3 == cnt[10:0] ? $signed(-32'shffbf) : $signed(_GEN_2019); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2021 = 11'h7e4 == cnt[10:0] ? $signed(-32'shffc4) : $signed(_GEN_2020); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2022 = 11'h7e5 == cnt[10:0] ? $signed(-32'shffc8) : $signed(_GEN_2021); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2023 = 11'h7e6 == cnt[10:0] ? $signed(-32'shffcc) : $signed(_GEN_2022); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2024 = 11'h7e7 == cnt[10:0] ? $signed(-32'shffd0) : $signed(_GEN_2023); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2025 = 11'h7e8 == cnt[10:0] ? $signed(-32'shffd4) : $signed(_GEN_2024); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2026 = 11'h7e9 == cnt[10:0] ? $signed(-32'shffd7) : $signed(_GEN_2025); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2027 = 11'h7ea == cnt[10:0] ? $signed(-32'shffdb) : $signed(_GEN_2026); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2028 = 11'h7eb == cnt[10:0] ? $signed(-32'shffde) : $signed(_GEN_2027); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2029 = 11'h7ec == cnt[10:0] ? $signed(-32'shffe1) : $signed(_GEN_2028); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2030 = 11'h7ed == cnt[10:0] ? $signed(-32'shffe4) : $signed(_GEN_2029); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2031 = 11'h7ee == cnt[10:0] ? $signed(-32'shffe7) : $signed(_GEN_2030); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2032 = 11'h7ef == cnt[10:0] ? $signed(-32'shffea) : $signed(_GEN_2031); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2033 = 11'h7f0 == cnt[10:0] ? $signed(-32'shffec) : $signed(_GEN_2032); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2034 = 11'h7f1 == cnt[10:0] ? $signed(-32'shffef) : $signed(_GEN_2033); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2035 = 11'h7f2 == cnt[10:0] ? $signed(-32'shfff1) : $signed(_GEN_2034); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2036 = 11'h7f3 == cnt[10:0] ? $signed(-32'shfff3) : $signed(_GEN_2035); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2037 = 11'h7f4 == cnt[10:0] ? $signed(-32'shfff5) : $signed(_GEN_2036); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2038 = 11'h7f5 == cnt[10:0] ? $signed(-32'shfff7) : $signed(_GEN_2037); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2039 = 11'h7f6 == cnt[10:0] ? $signed(-32'shfff8) : $signed(_GEN_2038); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2040 = 11'h7f7 == cnt[10:0] ? $signed(-32'shfffa) : $signed(_GEN_2039); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2041 = 11'h7f8 == cnt[10:0] ? $signed(-32'shfffb) : $signed(_GEN_2040); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2042 = 11'h7f9 == cnt[10:0] ? $signed(-32'shfffc) : $signed(_GEN_2041); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2043 = 11'h7fa == cnt[10:0] ? $signed(-32'shfffd) : $signed(_GEN_2042); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2044 = 11'h7fb == cnt[10:0] ? $signed(-32'shfffe) : $signed(_GEN_2043); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2045 = 11'h7fc == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_2044); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2046 = 11'h7fd == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_2045); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2047 = 11'h7fe == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_2046); // @[FFT.scala 34:12]
  wire [31:0] _GEN_2050 = 11'h1 == cnt[10:0] ? $signed(-32'sh65) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2051 = 11'h2 == cnt[10:0] ? $signed(-32'shc9) : $signed(_GEN_2050); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2052 = 11'h3 == cnt[10:0] ? $signed(-32'sh12e) : $signed(_GEN_2051); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2053 = 11'h4 == cnt[10:0] ? $signed(-32'sh192) : $signed(_GEN_2052); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2054 = 11'h5 == cnt[10:0] ? $signed(-32'sh1f7) : $signed(_GEN_2053); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2055 = 11'h6 == cnt[10:0] ? $signed(-32'sh25b) : $signed(_GEN_2054); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2056 = 11'h7 == cnt[10:0] ? $signed(-32'sh2c0) : $signed(_GEN_2055); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2057 = 11'h8 == cnt[10:0] ? $signed(-32'sh324) : $signed(_GEN_2056); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2058 = 11'h9 == cnt[10:0] ? $signed(-32'sh389) : $signed(_GEN_2057); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2059 = 11'ha == cnt[10:0] ? $signed(-32'sh3ed) : $signed(_GEN_2058); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2060 = 11'hb == cnt[10:0] ? $signed(-32'sh452) : $signed(_GEN_2059); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2061 = 11'hc == cnt[10:0] ? $signed(-32'sh4b6) : $signed(_GEN_2060); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2062 = 11'hd == cnt[10:0] ? $signed(-32'sh51b) : $signed(_GEN_2061); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2063 = 11'he == cnt[10:0] ? $signed(-32'sh57f) : $signed(_GEN_2062); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2064 = 11'hf == cnt[10:0] ? $signed(-32'sh5e4) : $signed(_GEN_2063); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2065 = 11'h10 == cnt[10:0] ? $signed(-32'sh648) : $signed(_GEN_2064); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2066 = 11'h11 == cnt[10:0] ? $signed(-32'sh6ad) : $signed(_GEN_2065); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2067 = 11'h12 == cnt[10:0] ? $signed(-32'sh711) : $signed(_GEN_2066); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2068 = 11'h13 == cnt[10:0] ? $signed(-32'sh776) : $signed(_GEN_2067); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2069 = 11'h14 == cnt[10:0] ? $signed(-32'sh7da) : $signed(_GEN_2068); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2070 = 11'h15 == cnt[10:0] ? $signed(-32'sh83f) : $signed(_GEN_2069); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2071 = 11'h16 == cnt[10:0] ? $signed(-32'sh8a3) : $signed(_GEN_2070); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2072 = 11'h17 == cnt[10:0] ? $signed(-32'sh908) : $signed(_GEN_2071); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2073 = 11'h18 == cnt[10:0] ? $signed(-32'sh96c) : $signed(_GEN_2072); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2074 = 11'h19 == cnt[10:0] ? $signed(-32'sh9d1) : $signed(_GEN_2073); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2075 = 11'h1a == cnt[10:0] ? $signed(-32'sha35) : $signed(_GEN_2074); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2076 = 11'h1b == cnt[10:0] ? $signed(-32'sha9a) : $signed(_GEN_2075); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2077 = 11'h1c == cnt[10:0] ? $signed(-32'shafe) : $signed(_GEN_2076); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2078 = 11'h1d == cnt[10:0] ? $signed(-32'shb62) : $signed(_GEN_2077); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2079 = 11'h1e == cnt[10:0] ? $signed(-32'shbc7) : $signed(_GEN_2078); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2080 = 11'h1f == cnt[10:0] ? $signed(-32'shc2b) : $signed(_GEN_2079); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2081 = 11'h20 == cnt[10:0] ? $signed(-32'shc90) : $signed(_GEN_2080); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2082 = 11'h21 == cnt[10:0] ? $signed(-32'shcf4) : $signed(_GEN_2081); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2083 = 11'h22 == cnt[10:0] ? $signed(-32'shd59) : $signed(_GEN_2082); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2084 = 11'h23 == cnt[10:0] ? $signed(-32'shdbd) : $signed(_GEN_2083); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2085 = 11'h24 == cnt[10:0] ? $signed(-32'she21) : $signed(_GEN_2084); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2086 = 11'h25 == cnt[10:0] ? $signed(-32'she86) : $signed(_GEN_2085); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2087 = 11'h26 == cnt[10:0] ? $signed(-32'sheea) : $signed(_GEN_2086); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2088 = 11'h27 == cnt[10:0] ? $signed(-32'shf4e) : $signed(_GEN_2087); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2089 = 11'h28 == cnt[10:0] ? $signed(-32'shfb3) : $signed(_GEN_2088); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2090 = 11'h29 == cnt[10:0] ? $signed(-32'sh1017) : $signed(_GEN_2089); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2091 = 11'h2a == cnt[10:0] ? $signed(-32'sh107b) : $signed(_GEN_2090); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2092 = 11'h2b == cnt[10:0] ? $signed(-32'sh10e0) : $signed(_GEN_2091); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2093 = 11'h2c == cnt[10:0] ? $signed(-32'sh1144) : $signed(_GEN_2092); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2094 = 11'h2d == cnt[10:0] ? $signed(-32'sh11a8) : $signed(_GEN_2093); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2095 = 11'h2e == cnt[10:0] ? $signed(-32'sh120d) : $signed(_GEN_2094); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2096 = 11'h2f == cnt[10:0] ? $signed(-32'sh1271) : $signed(_GEN_2095); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2097 = 11'h30 == cnt[10:0] ? $signed(-32'sh12d5) : $signed(_GEN_2096); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2098 = 11'h31 == cnt[10:0] ? $signed(-32'sh1339) : $signed(_GEN_2097); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2099 = 11'h32 == cnt[10:0] ? $signed(-32'sh139e) : $signed(_GEN_2098); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2100 = 11'h33 == cnt[10:0] ? $signed(-32'sh1402) : $signed(_GEN_2099); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2101 = 11'h34 == cnt[10:0] ? $signed(-32'sh1466) : $signed(_GEN_2100); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2102 = 11'h35 == cnt[10:0] ? $signed(-32'sh14ca) : $signed(_GEN_2101); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2103 = 11'h36 == cnt[10:0] ? $signed(-32'sh152e) : $signed(_GEN_2102); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2104 = 11'h37 == cnt[10:0] ? $signed(-32'sh1593) : $signed(_GEN_2103); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2105 = 11'h38 == cnt[10:0] ? $signed(-32'sh15f7) : $signed(_GEN_2104); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2106 = 11'h39 == cnt[10:0] ? $signed(-32'sh165b) : $signed(_GEN_2105); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2107 = 11'h3a == cnt[10:0] ? $signed(-32'sh16bf) : $signed(_GEN_2106); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2108 = 11'h3b == cnt[10:0] ? $signed(-32'sh1723) : $signed(_GEN_2107); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2109 = 11'h3c == cnt[10:0] ? $signed(-32'sh1787) : $signed(_GEN_2108); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2110 = 11'h3d == cnt[10:0] ? $signed(-32'sh17eb) : $signed(_GEN_2109); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2111 = 11'h3e == cnt[10:0] ? $signed(-32'sh1850) : $signed(_GEN_2110); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2112 = 11'h3f == cnt[10:0] ? $signed(-32'sh18b4) : $signed(_GEN_2111); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2113 = 11'h40 == cnt[10:0] ? $signed(-32'sh1918) : $signed(_GEN_2112); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2114 = 11'h41 == cnt[10:0] ? $signed(-32'sh197c) : $signed(_GEN_2113); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2115 = 11'h42 == cnt[10:0] ? $signed(-32'sh19e0) : $signed(_GEN_2114); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2116 = 11'h43 == cnt[10:0] ? $signed(-32'sh1a44) : $signed(_GEN_2115); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2117 = 11'h44 == cnt[10:0] ? $signed(-32'sh1aa8) : $signed(_GEN_2116); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2118 = 11'h45 == cnt[10:0] ? $signed(-32'sh1b0c) : $signed(_GEN_2117); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2119 = 11'h46 == cnt[10:0] ? $signed(-32'sh1b70) : $signed(_GEN_2118); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2120 = 11'h47 == cnt[10:0] ? $signed(-32'sh1bd4) : $signed(_GEN_2119); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2121 = 11'h48 == cnt[10:0] ? $signed(-32'sh1c38) : $signed(_GEN_2120); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2122 = 11'h49 == cnt[10:0] ? $signed(-32'sh1c9b) : $signed(_GEN_2121); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2123 = 11'h4a == cnt[10:0] ? $signed(-32'sh1cff) : $signed(_GEN_2122); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2124 = 11'h4b == cnt[10:0] ? $signed(-32'sh1d63) : $signed(_GEN_2123); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2125 = 11'h4c == cnt[10:0] ? $signed(-32'sh1dc7) : $signed(_GEN_2124); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2126 = 11'h4d == cnt[10:0] ? $signed(-32'sh1e2b) : $signed(_GEN_2125); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2127 = 11'h4e == cnt[10:0] ? $signed(-32'sh1e8f) : $signed(_GEN_2126); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2128 = 11'h4f == cnt[10:0] ? $signed(-32'sh1ef3) : $signed(_GEN_2127); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2129 = 11'h50 == cnt[10:0] ? $signed(-32'sh1f56) : $signed(_GEN_2128); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2130 = 11'h51 == cnt[10:0] ? $signed(-32'sh1fba) : $signed(_GEN_2129); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2131 = 11'h52 == cnt[10:0] ? $signed(-32'sh201e) : $signed(_GEN_2130); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2132 = 11'h53 == cnt[10:0] ? $signed(-32'sh2082) : $signed(_GEN_2131); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2133 = 11'h54 == cnt[10:0] ? $signed(-32'sh20e5) : $signed(_GEN_2132); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2134 = 11'h55 == cnt[10:0] ? $signed(-32'sh2149) : $signed(_GEN_2133); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2135 = 11'h56 == cnt[10:0] ? $signed(-32'sh21ad) : $signed(_GEN_2134); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2136 = 11'h57 == cnt[10:0] ? $signed(-32'sh2210) : $signed(_GEN_2135); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2137 = 11'h58 == cnt[10:0] ? $signed(-32'sh2274) : $signed(_GEN_2136); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2138 = 11'h59 == cnt[10:0] ? $signed(-32'sh22d7) : $signed(_GEN_2137); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2139 = 11'h5a == cnt[10:0] ? $signed(-32'sh233b) : $signed(_GEN_2138); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2140 = 11'h5b == cnt[10:0] ? $signed(-32'sh239f) : $signed(_GEN_2139); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2141 = 11'h5c == cnt[10:0] ? $signed(-32'sh2402) : $signed(_GEN_2140); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2142 = 11'h5d == cnt[10:0] ? $signed(-32'sh2466) : $signed(_GEN_2141); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2143 = 11'h5e == cnt[10:0] ? $signed(-32'sh24c9) : $signed(_GEN_2142); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2144 = 11'h5f == cnt[10:0] ? $signed(-32'sh252d) : $signed(_GEN_2143); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2145 = 11'h60 == cnt[10:0] ? $signed(-32'sh2590) : $signed(_GEN_2144); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2146 = 11'h61 == cnt[10:0] ? $signed(-32'sh25f4) : $signed(_GEN_2145); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2147 = 11'h62 == cnt[10:0] ? $signed(-32'sh2657) : $signed(_GEN_2146); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2148 = 11'h63 == cnt[10:0] ? $signed(-32'sh26ba) : $signed(_GEN_2147); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2149 = 11'h64 == cnt[10:0] ? $signed(-32'sh271e) : $signed(_GEN_2148); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2150 = 11'h65 == cnt[10:0] ? $signed(-32'sh2781) : $signed(_GEN_2149); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2151 = 11'h66 == cnt[10:0] ? $signed(-32'sh27e4) : $signed(_GEN_2150); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2152 = 11'h67 == cnt[10:0] ? $signed(-32'sh2848) : $signed(_GEN_2151); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2153 = 11'h68 == cnt[10:0] ? $signed(-32'sh28ab) : $signed(_GEN_2152); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2154 = 11'h69 == cnt[10:0] ? $signed(-32'sh290e) : $signed(_GEN_2153); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2155 = 11'h6a == cnt[10:0] ? $signed(-32'sh2971) : $signed(_GEN_2154); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2156 = 11'h6b == cnt[10:0] ? $signed(-32'sh29d5) : $signed(_GEN_2155); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2157 = 11'h6c == cnt[10:0] ? $signed(-32'sh2a38) : $signed(_GEN_2156); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2158 = 11'h6d == cnt[10:0] ? $signed(-32'sh2a9b) : $signed(_GEN_2157); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2159 = 11'h6e == cnt[10:0] ? $signed(-32'sh2afe) : $signed(_GEN_2158); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2160 = 11'h6f == cnt[10:0] ? $signed(-32'sh2b61) : $signed(_GEN_2159); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2161 = 11'h70 == cnt[10:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2160); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2162 = 11'h71 == cnt[10:0] ? $signed(-32'sh2c27) : $signed(_GEN_2161); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2163 = 11'h72 == cnt[10:0] ? $signed(-32'sh2c8a) : $signed(_GEN_2162); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2164 = 11'h73 == cnt[10:0] ? $signed(-32'sh2ced) : $signed(_GEN_2163); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2165 = 11'h74 == cnt[10:0] ? $signed(-32'sh2d50) : $signed(_GEN_2164); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2166 = 11'h75 == cnt[10:0] ? $signed(-32'sh2db3) : $signed(_GEN_2165); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2167 = 11'h76 == cnt[10:0] ? $signed(-32'sh2e16) : $signed(_GEN_2166); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2168 = 11'h77 == cnt[10:0] ? $signed(-32'sh2e79) : $signed(_GEN_2167); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2169 = 11'h78 == cnt[10:0] ? $signed(-32'sh2edc) : $signed(_GEN_2168); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2170 = 11'h79 == cnt[10:0] ? $signed(-32'sh2f3f) : $signed(_GEN_2169); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2171 = 11'h7a == cnt[10:0] ? $signed(-32'sh2fa1) : $signed(_GEN_2170); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2172 = 11'h7b == cnt[10:0] ? $signed(-32'sh3004) : $signed(_GEN_2171); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2173 = 11'h7c == cnt[10:0] ? $signed(-32'sh3067) : $signed(_GEN_2172); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2174 = 11'h7d == cnt[10:0] ? $signed(-32'sh30ca) : $signed(_GEN_2173); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2175 = 11'h7e == cnt[10:0] ? $signed(-32'sh312c) : $signed(_GEN_2174); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2176 = 11'h7f == cnt[10:0] ? $signed(-32'sh318f) : $signed(_GEN_2175); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2177 = 11'h80 == cnt[10:0] ? $signed(-32'sh31f1) : $signed(_GEN_2176); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2178 = 11'h81 == cnt[10:0] ? $signed(-32'sh3254) : $signed(_GEN_2177); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2179 = 11'h82 == cnt[10:0] ? $signed(-32'sh32b7) : $signed(_GEN_2178); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2180 = 11'h83 == cnt[10:0] ? $signed(-32'sh3319) : $signed(_GEN_2179); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2181 = 11'h84 == cnt[10:0] ? $signed(-32'sh337c) : $signed(_GEN_2180); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2182 = 11'h85 == cnt[10:0] ? $signed(-32'sh33de) : $signed(_GEN_2181); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2183 = 11'h86 == cnt[10:0] ? $signed(-32'sh3440) : $signed(_GEN_2182); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2184 = 11'h87 == cnt[10:0] ? $signed(-32'sh34a3) : $signed(_GEN_2183); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2185 = 11'h88 == cnt[10:0] ? $signed(-32'sh3505) : $signed(_GEN_2184); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2186 = 11'h89 == cnt[10:0] ? $signed(-32'sh3568) : $signed(_GEN_2185); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2187 = 11'h8a == cnt[10:0] ? $signed(-32'sh35ca) : $signed(_GEN_2186); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2188 = 11'h8b == cnt[10:0] ? $signed(-32'sh362c) : $signed(_GEN_2187); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2189 = 11'h8c == cnt[10:0] ? $signed(-32'sh368e) : $signed(_GEN_2188); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2190 = 11'h8d == cnt[10:0] ? $signed(-32'sh36f1) : $signed(_GEN_2189); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2191 = 11'h8e == cnt[10:0] ? $signed(-32'sh3753) : $signed(_GEN_2190); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2192 = 11'h8f == cnt[10:0] ? $signed(-32'sh37b5) : $signed(_GEN_2191); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2193 = 11'h90 == cnt[10:0] ? $signed(-32'sh3817) : $signed(_GEN_2192); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2194 = 11'h91 == cnt[10:0] ? $signed(-32'sh3879) : $signed(_GEN_2193); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2195 = 11'h92 == cnt[10:0] ? $signed(-32'sh38db) : $signed(_GEN_2194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2196 = 11'h93 == cnt[10:0] ? $signed(-32'sh393d) : $signed(_GEN_2195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2197 = 11'h94 == cnt[10:0] ? $signed(-32'sh399f) : $signed(_GEN_2196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2198 = 11'h95 == cnt[10:0] ? $signed(-32'sh3a01) : $signed(_GEN_2197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2199 = 11'h96 == cnt[10:0] ? $signed(-32'sh3a63) : $signed(_GEN_2198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2200 = 11'h97 == cnt[10:0] ? $signed(-32'sh3ac5) : $signed(_GEN_2199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2201 = 11'h98 == cnt[10:0] ? $signed(-32'sh3b27) : $signed(_GEN_2200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2202 = 11'h99 == cnt[10:0] ? $signed(-32'sh3b88) : $signed(_GEN_2201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2203 = 11'h9a == cnt[10:0] ? $signed(-32'sh3bea) : $signed(_GEN_2202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2204 = 11'h9b == cnt[10:0] ? $signed(-32'sh3c4c) : $signed(_GEN_2203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2205 = 11'h9c == cnt[10:0] ? $signed(-32'sh3cae) : $signed(_GEN_2204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2206 = 11'h9d == cnt[10:0] ? $signed(-32'sh3d0f) : $signed(_GEN_2205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2207 = 11'h9e == cnt[10:0] ? $signed(-32'sh3d71) : $signed(_GEN_2206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2208 = 11'h9f == cnt[10:0] ? $signed(-32'sh3dd2) : $signed(_GEN_2207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2209 = 11'ha0 == cnt[10:0] ? $signed(-32'sh3e34) : $signed(_GEN_2208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2210 = 11'ha1 == cnt[10:0] ? $signed(-32'sh3e95) : $signed(_GEN_2209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2211 = 11'ha2 == cnt[10:0] ? $signed(-32'sh3ef7) : $signed(_GEN_2210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2212 = 11'ha3 == cnt[10:0] ? $signed(-32'sh3f58) : $signed(_GEN_2211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2213 = 11'ha4 == cnt[10:0] ? $signed(-32'sh3fba) : $signed(_GEN_2212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2214 = 11'ha5 == cnt[10:0] ? $signed(-32'sh401b) : $signed(_GEN_2213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2215 = 11'ha6 == cnt[10:0] ? $signed(-32'sh407c) : $signed(_GEN_2214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2216 = 11'ha7 == cnt[10:0] ? $signed(-32'sh40de) : $signed(_GEN_2215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2217 = 11'ha8 == cnt[10:0] ? $signed(-32'sh413f) : $signed(_GEN_2216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2218 = 11'ha9 == cnt[10:0] ? $signed(-32'sh41a0) : $signed(_GEN_2217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2219 = 11'haa == cnt[10:0] ? $signed(-32'sh4201) : $signed(_GEN_2218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2220 = 11'hab == cnt[10:0] ? $signed(-32'sh4262) : $signed(_GEN_2219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2221 = 11'hac == cnt[10:0] ? $signed(-32'sh42c3) : $signed(_GEN_2220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2222 = 11'had == cnt[10:0] ? $signed(-32'sh4324) : $signed(_GEN_2221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2223 = 11'hae == cnt[10:0] ? $signed(-32'sh4385) : $signed(_GEN_2222); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2224 = 11'haf == cnt[10:0] ? $signed(-32'sh43e6) : $signed(_GEN_2223); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2225 = 11'hb0 == cnt[10:0] ? $signed(-32'sh4447) : $signed(_GEN_2224); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2226 = 11'hb1 == cnt[10:0] ? $signed(-32'sh44a8) : $signed(_GEN_2225); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2227 = 11'hb2 == cnt[10:0] ? $signed(-32'sh4509) : $signed(_GEN_2226); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2228 = 11'hb3 == cnt[10:0] ? $signed(-32'sh456a) : $signed(_GEN_2227); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2229 = 11'hb4 == cnt[10:0] ? $signed(-32'sh45cb) : $signed(_GEN_2228); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2230 = 11'hb5 == cnt[10:0] ? $signed(-32'sh462b) : $signed(_GEN_2229); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2231 = 11'hb6 == cnt[10:0] ? $signed(-32'sh468c) : $signed(_GEN_2230); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2232 = 11'hb7 == cnt[10:0] ? $signed(-32'sh46ec) : $signed(_GEN_2231); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2233 = 11'hb8 == cnt[10:0] ? $signed(-32'sh474d) : $signed(_GEN_2232); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2234 = 11'hb9 == cnt[10:0] ? $signed(-32'sh47ae) : $signed(_GEN_2233); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2235 = 11'hba == cnt[10:0] ? $signed(-32'sh480e) : $signed(_GEN_2234); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2236 = 11'hbb == cnt[10:0] ? $signed(-32'sh486f) : $signed(_GEN_2235); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2237 = 11'hbc == cnt[10:0] ? $signed(-32'sh48cf) : $signed(_GEN_2236); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2238 = 11'hbd == cnt[10:0] ? $signed(-32'sh492f) : $signed(_GEN_2237); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2239 = 11'hbe == cnt[10:0] ? $signed(-32'sh4990) : $signed(_GEN_2238); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2240 = 11'hbf == cnt[10:0] ? $signed(-32'sh49f0) : $signed(_GEN_2239); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2241 = 11'hc0 == cnt[10:0] ? $signed(-32'sh4a50) : $signed(_GEN_2240); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2242 = 11'hc1 == cnt[10:0] ? $signed(-32'sh4ab0) : $signed(_GEN_2241); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2243 = 11'hc2 == cnt[10:0] ? $signed(-32'sh4b10) : $signed(_GEN_2242); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2244 = 11'hc3 == cnt[10:0] ? $signed(-32'sh4b71) : $signed(_GEN_2243); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2245 = 11'hc4 == cnt[10:0] ? $signed(-32'sh4bd1) : $signed(_GEN_2244); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2246 = 11'hc5 == cnt[10:0] ? $signed(-32'sh4c31) : $signed(_GEN_2245); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2247 = 11'hc6 == cnt[10:0] ? $signed(-32'sh4c90) : $signed(_GEN_2246); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2248 = 11'hc7 == cnt[10:0] ? $signed(-32'sh4cf0) : $signed(_GEN_2247); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2249 = 11'hc8 == cnt[10:0] ? $signed(-32'sh4d50) : $signed(_GEN_2248); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2250 = 11'hc9 == cnt[10:0] ? $signed(-32'sh4db0) : $signed(_GEN_2249); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2251 = 11'hca == cnt[10:0] ? $signed(-32'sh4e10) : $signed(_GEN_2250); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2252 = 11'hcb == cnt[10:0] ? $signed(-32'sh4e70) : $signed(_GEN_2251); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2253 = 11'hcc == cnt[10:0] ? $signed(-32'sh4ecf) : $signed(_GEN_2252); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2254 = 11'hcd == cnt[10:0] ? $signed(-32'sh4f2f) : $signed(_GEN_2253); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2255 = 11'hce == cnt[10:0] ? $signed(-32'sh4f8e) : $signed(_GEN_2254); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2256 = 11'hcf == cnt[10:0] ? $signed(-32'sh4fee) : $signed(_GEN_2255); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2257 = 11'hd0 == cnt[10:0] ? $signed(-32'sh504d) : $signed(_GEN_2256); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2258 = 11'hd1 == cnt[10:0] ? $signed(-32'sh50ad) : $signed(_GEN_2257); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2259 = 11'hd2 == cnt[10:0] ? $signed(-32'sh510c) : $signed(_GEN_2258); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2260 = 11'hd3 == cnt[10:0] ? $signed(-32'sh516c) : $signed(_GEN_2259); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2261 = 11'hd4 == cnt[10:0] ? $signed(-32'sh51cb) : $signed(_GEN_2260); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2262 = 11'hd5 == cnt[10:0] ? $signed(-32'sh522a) : $signed(_GEN_2261); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2263 = 11'hd6 == cnt[10:0] ? $signed(-32'sh5289) : $signed(_GEN_2262); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2264 = 11'hd7 == cnt[10:0] ? $signed(-32'sh52e8) : $signed(_GEN_2263); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2265 = 11'hd8 == cnt[10:0] ? $signed(-32'sh5348) : $signed(_GEN_2264); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2266 = 11'hd9 == cnt[10:0] ? $signed(-32'sh53a7) : $signed(_GEN_2265); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2267 = 11'hda == cnt[10:0] ? $signed(-32'sh5406) : $signed(_GEN_2266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2268 = 11'hdb == cnt[10:0] ? $signed(-32'sh5464) : $signed(_GEN_2267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2269 = 11'hdc == cnt[10:0] ? $signed(-32'sh54c3) : $signed(_GEN_2268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2270 = 11'hdd == cnt[10:0] ? $signed(-32'sh5522) : $signed(_GEN_2269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2271 = 11'hde == cnt[10:0] ? $signed(-32'sh5581) : $signed(_GEN_2270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2272 = 11'hdf == cnt[10:0] ? $signed(-32'sh55e0) : $signed(_GEN_2271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2273 = 11'he0 == cnt[10:0] ? $signed(-32'sh563e) : $signed(_GEN_2272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2274 = 11'he1 == cnt[10:0] ? $signed(-32'sh569d) : $signed(_GEN_2273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2275 = 11'he2 == cnt[10:0] ? $signed(-32'sh56fc) : $signed(_GEN_2274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2276 = 11'he3 == cnt[10:0] ? $signed(-32'sh575a) : $signed(_GEN_2275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2277 = 11'he4 == cnt[10:0] ? $signed(-32'sh57b9) : $signed(_GEN_2276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2278 = 11'he5 == cnt[10:0] ? $signed(-32'sh5817) : $signed(_GEN_2277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2279 = 11'he6 == cnt[10:0] ? $signed(-32'sh5875) : $signed(_GEN_2278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2280 = 11'he7 == cnt[10:0] ? $signed(-32'sh58d4) : $signed(_GEN_2279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2281 = 11'he8 == cnt[10:0] ? $signed(-32'sh5932) : $signed(_GEN_2280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2282 = 11'he9 == cnt[10:0] ? $signed(-32'sh5990) : $signed(_GEN_2281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2283 = 11'hea == cnt[10:0] ? $signed(-32'sh59ee) : $signed(_GEN_2282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2284 = 11'heb == cnt[10:0] ? $signed(-32'sh5a4c) : $signed(_GEN_2283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2285 = 11'hec == cnt[10:0] ? $signed(-32'sh5aaa) : $signed(_GEN_2284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2286 = 11'hed == cnt[10:0] ? $signed(-32'sh5b08) : $signed(_GEN_2285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2287 = 11'hee == cnt[10:0] ? $signed(-32'sh5b66) : $signed(_GEN_2286); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2288 = 11'hef == cnt[10:0] ? $signed(-32'sh5bc4) : $signed(_GEN_2287); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2289 = 11'hf0 == cnt[10:0] ? $signed(-32'sh5c22) : $signed(_GEN_2288); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2290 = 11'hf1 == cnt[10:0] ? $signed(-32'sh5c80) : $signed(_GEN_2289); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2291 = 11'hf2 == cnt[10:0] ? $signed(-32'sh5cde) : $signed(_GEN_2290); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2292 = 11'hf3 == cnt[10:0] ? $signed(-32'sh5d3b) : $signed(_GEN_2291); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2293 = 11'hf4 == cnt[10:0] ? $signed(-32'sh5d99) : $signed(_GEN_2292); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2294 = 11'hf5 == cnt[10:0] ? $signed(-32'sh5df6) : $signed(_GEN_2293); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2295 = 11'hf6 == cnt[10:0] ? $signed(-32'sh5e54) : $signed(_GEN_2294); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2296 = 11'hf7 == cnt[10:0] ? $signed(-32'sh5eb1) : $signed(_GEN_2295); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2297 = 11'hf8 == cnt[10:0] ? $signed(-32'sh5f0f) : $signed(_GEN_2296); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2298 = 11'hf9 == cnt[10:0] ? $signed(-32'sh5f6c) : $signed(_GEN_2297); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2299 = 11'hfa == cnt[10:0] ? $signed(-32'sh5fc9) : $signed(_GEN_2298); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2300 = 11'hfb == cnt[10:0] ? $signed(-32'sh6026) : $signed(_GEN_2299); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2301 = 11'hfc == cnt[10:0] ? $signed(-32'sh6084) : $signed(_GEN_2300); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2302 = 11'hfd == cnt[10:0] ? $signed(-32'sh60e1) : $signed(_GEN_2301); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2303 = 11'hfe == cnt[10:0] ? $signed(-32'sh613e) : $signed(_GEN_2302); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2304 = 11'hff == cnt[10:0] ? $signed(-32'sh619b) : $signed(_GEN_2303); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2305 = 11'h100 == cnt[10:0] ? $signed(-32'sh61f8) : $signed(_GEN_2304); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2306 = 11'h101 == cnt[10:0] ? $signed(-32'sh6254) : $signed(_GEN_2305); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2307 = 11'h102 == cnt[10:0] ? $signed(-32'sh62b1) : $signed(_GEN_2306); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2308 = 11'h103 == cnt[10:0] ? $signed(-32'sh630e) : $signed(_GEN_2307); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2309 = 11'h104 == cnt[10:0] ? $signed(-32'sh636b) : $signed(_GEN_2308); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2310 = 11'h105 == cnt[10:0] ? $signed(-32'sh63c7) : $signed(_GEN_2309); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2311 = 11'h106 == cnt[10:0] ? $signed(-32'sh6424) : $signed(_GEN_2310); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2312 = 11'h107 == cnt[10:0] ? $signed(-32'sh6480) : $signed(_GEN_2311); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2313 = 11'h108 == cnt[10:0] ? $signed(-32'sh64dd) : $signed(_GEN_2312); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2314 = 11'h109 == cnt[10:0] ? $signed(-32'sh6539) : $signed(_GEN_2313); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2315 = 11'h10a == cnt[10:0] ? $signed(-32'sh6595) : $signed(_GEN_2314); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2316 = 11'h10b == cnt[10:0] ? $signed(-32'sh65f2) : $signed(_GEN_2315); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2317 = 11'h10c == cnt[10:0] ? $signed(-32'sh664e) : $signed(_GEN_2316); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2318 = 11'h10d == cnt[10:0] ? $signed(-32'sh66aa) : $signed(_GEN_2317); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2319 = 11'h10e == cnt[10:0] ? $signed(-32'sh6706) : $signed(_GEN_2318); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2320 = 11'h10f == cnt[10:0] ? $signed(-32'sh6762) : $signed(_GEN_2319); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2321 = 11'h110 == cnt[10:0] ? $signed(-32'sh67be) : $signed(_GEN_2320); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2322 = 11'h111 == cnt[10:0] ? $signed(-32'sh681a) : $signed(_GEN_2321); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2323 = 11'h112 == cnt[10:0] ? $signed(-32'sh6876) : $signed(_GEN_2322); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2324 = 11'h113 == cnt[10:0] ? $signed(-32'sh68d1) : $signed(_GEN_2323); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2325 = 11'h114 == cnt[10:0] ? $signed(-32'sh692d) : $signed(_GEN_2324); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2326 = 11'h115 == cnt[10:0] ? $signed(-32'sh6989) : $signed(_GEN_2325); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2327 = 11'h116 == cnt[10:0] ? $signed(-32'sh69e4) : $signed(_GEN_2326); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2328 = 11'h117 == cnt[10:0] ? $signed(-32'sh6a40) : $signed(_GEN_2327); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2329 = 11'h118 == cnt[10:0] ? $signed(-32'sh6a9b) : $signed(_GEN_2328); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2330 = 11'h119 == cnt[10:0] ? $signed(-32'sh6af6) : $signed(_GEN_2329); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2331 = 11'h11a == cnt[10:0] ? $signed(-32'sh6b52) : $signed(_GEN_2330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2332 = 11'h11b == cnt[10:0] ? $signed(-32'sh6bad) : $signed(_GEN_2331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2333 = 11'h11c == cnt[10:0] ? $signed(-32'sh6c08) : $signed(_GEN_2332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2334 = 11'h11d == cnt[10:0] ? $signed(-32'sh6c63) : $signed(_GEN_2333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2335 = 11'h11e == cnt[10:0] ? $signed(-32'sh6cbe) : $signed(_GEN_2334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2336 = 11'h11f == cnt[10:0] ? $signed(-32'sh6d19) : $signed(_GEN_2335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2337 = 11'h120 == cnt[10:0] ? $signed(-32'sh6d74) : $signed(_GEN_2336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2338 = 11'h121 == cnt[10:0] ? $signed(-32'sh6dcf) : $signed(_GEN_2337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2339 = 11'h122 == cnt[10:0] ? $signed(-32'sh6e2a) : $signed(_GEN_2338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2340 = 11'h123 == cnt[10:0] ? $signed(-32'sh6e85) : $signed(_GEN_2339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2341 = 11'h124 == cnt[10:0] ? $signed(-32'sh6edf) : $signed(_GEN_2340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2342 = 11'h125 == cnt[10:0] ? $signed(-32'sh6f3a) : $signed(_GEN_2341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2343 = 11'h126 == cnt[10:0] ? $signed(-32'sh6f94) : $signed(_GEN_2342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2344 = 11'h127 == cnt[10:0] ? $signed(-32'sh6fef) : $signed(_GEN_2343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2345 = 11'h128 == cnt[10:0] ? $signed(-32'sh7049) : $signed(_GEN_2344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2346 = 11'h129 == cnt[10:0] ? $signed(-32'sh70a3) : $signed(_GEN_2345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2347 = 11'h12a == cnt[10:0] ? $signed(-32'sh70fe) : $signed(_GEN_2346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2348 = 11'h12b == cnt[10:0] ? $signed(-32'sh7158) : $signed(_GEN_2347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2349 = 11'h12c == cnt[10:0] ? $signed(-32'sh71b2) : $signed(_GEN_2348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2350 = 11'h12d == cnt[10:0] ? $signed(-32'sh720c) : $signed(_GEN_2349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2351 = 11'h12e == cnt[10:0] ? $signed(-32'sh7266) : $signed(_GEN_2350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2352 = 11'h12f == cnt[10:0] ? $signed(-32'sh72c0) : $signed(_GEN_2351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2353 = 11'h130 == cnt[10:0] ? $signed(-32'sh731a) : $signed(_GEN_2352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2354 = 11'h131 == cnt[10:0] ? $signed(-32'sh7373) : $signed(_GEN_2353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2355 = 11'h132 == cnt[10:0] ? $signed(-32'sh73cd) : $signed(_GEN_2354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2356 = 11'h133 == cnt[10:0] ? $signed(-32'sh7427) : $signed(_GEN_2355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2357 = 11'h134 == cnt[10:0] ? $signed(-32'sh7480) : $signed(_GEN_2356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2358 = 11'h135 == cnt[10:0] ? $signed(-32'sh74da) : $signed(_GEN_2357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2359 = 11'h136 == cnt[10:0] ? $signed(-32'sh7533) : $signed(_GEN_2358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2360 = 11'h137 == cnt[10:0] ? $signed(-32'sh758d) : $signed(_GEN_2359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2361 = 11'h138 == cnt[10:0] ? $signed(-32'sh75e6) : $signed(_GEN_2360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2362 = 11'h139 == cnt[10:0] ? $signed(-32'sh763f) : $signed(_GEN_2361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2363 = 11'h13a == cnt[10:0] ? $signed(-32'sh7698) : $signed(_GEN_2362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2364 = 11'h13b == cnt[10:0] ? $signed(-32'sh76f1) : $signed(_GEN_2363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2365 = 11'h13c == cnt[10:0] ? $signed(-32'sh774a) : $signed(_GEN_2364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2366 = 11'h13d == cnt[10:0] ? $signed(-32'sh77a3) : $signed(_GEN_2365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2367 = 11'h13e == cnt[10:0] ? $signed(-32'sh77fc) : $signed(_GEN_2366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2368 = 11'h13f == cnt[10:0] ? $signed(-32'sh7855) : $signed(_GEN_2367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2369 = 11'h140 == cnt[10:0] ? $signed(-32'sh78ad) : $signed(_GEN_2368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2370 = 11'h141 == cnt[10:0] ? $signed(-32'sh7906) : $signed(_GEN_2369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2371 = 11'h142 == cnt[10:0] ? $signed(-32'sh795f) : $signed(_GEN_2370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2372 = 11'h143 == cnt[10:0] ? $signed(-32'sh79b7) : $signed(_GEN_2371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2373 = 11'h144 == cnt[10:0] ? $signed(-32'sh7a10) : $signed(_GEN_2372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2374 = 11'h145 == cnt[10:0] ? $signed(-32'sh7a68) : $signed(_GEN_2373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2375 = 11'h146 == cnt[10:0] ? $signed(-32'sh7ac0) : $signed(_GEN_2374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2376 = 11'h147 == cnt[10:0] ? $signed(-32'sh7b18) : $signed(_GEN_2375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2377 = 11'h148 == cnt[10:0] ? $signed(-32'sh7b70) : $signed(_GEN_2376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2378 = 11'h149 == cnt[10:0] ? $signed(-32'sh7bc8) : $signed(_GEN_2377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2379 = 11'h14a == cnt[10:0] ? $signed(-32'sh7c20) : $signed(_GEN_2378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2380 = 11'h14b == cnt[10:0] ? $signed(-32'sh7c78) : $signed(_GEN_2379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2381 = 11'h14c == cnt[10:0] ? $signed(-32'sh7cd0) : $signed(_GEN_2380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2382 = 11'h14d == cnt[10:0] ? $signed(-32'sh7d28) : $signed(_GEN_2381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2383 = 11'h14e == cnt[10:0] ? $signed(-32'sh7d7f) : $signed(_GEN_2382); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2384 = 11'h14f == cnt[10:0] ? $signed(-32'sh7dd7) : $signed(_GEN_2383); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2385 = 11'h150 == cnt[10:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2384); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2386 = 11'h151 == cnt[10:0] ? $signed(-32'sh7e86) : $signed(_GEN_2385); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2387 = 11'h152 == cnt[10:0] ? $signed(-32'sh7edd) : $signed(_GEN_2386); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2388 = 11'h153 == cnt[10:0] ? $signed(-32'sh7f35) : $signed(_GEN_2387); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2389 = 11'h154 == cnt[10:0] ? $signed(-32'sh7f8c) : $signed(_GEN_2388); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2390 = 11'h155 == cnt[10:0] ? $signed(-32'sh7fe3) : $signed(_GEN_2389); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2391 = 11'h156 == cnt[10:0] ? $signed(-32'sh803a) : $signed(_GEN_2390); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2392 = 11'h157 == cnt[10:0] ? $signed(-32'sh8091) : $signed(_GEN_2391); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2393 = 11'h158 == cnt[10:0] ? $signed(-32'sh80e8) : $signed(_GEN_2392); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2394 = 11'h159 == cnt[10:0] ? $signed(-32'sh813f) : $signed(_GEN_2393); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2395 = 11'h15a == cnt[10:0] ? $signed(-32'sh8195) : $signed(_GEN_2394); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2396 = 11'h15b == cnt[10:0] ? $signed(-32'sh81ec) : $signed(_GEN_2395); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2397 = 11'h15c == cnt[10:0] ? $signed(-32'sh8243) : $signed(_GEN_2396); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2398 = 11'h15d == cnt[10:0] ? $signed(-32'sh8299) : $signed(_GEN_2397); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2399 = 11'h15e == cnt[10:0] ? $signed(-32'sh82f0) : $signed(_GEN_2398); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2400 = 11'h15f == cnt[10:0] ? $signed(-32'sh8346) : $signed(_GEN_2399); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2401 = 11'h160 == cnt[10:0] ? $signed(-32'sh839c) : $signed(_GEN_2400); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2402 = 11'h161 == cnt[10:0] ? $signed(-32'sh83f2) : $signed(_GEN_2401); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2403 = 11'h162 == cnt[10:0] ? $signed(-32'sh8449) : $signed(_GEN_2402); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2404 = 11'h163 == cnt[10:0] ? $signed(-32'sh849f) : $signed(_GEN_2403); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2405 = 11'h164 == cnt[10:0] ? $signed(-32'sh84f5) : $signed(_GEN_2404); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2406 = 11'h165 == cnt[10:0] ? $signed(-32'sh854a) : $signed(_GEN_2405); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2407 = 11'h166 == cnt[10:0] ? $signed(-32'sh85a0) : $signed(_GEN_2406); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2408 = 11'h167 == cnt[10:0] ? $signed(-32'sh85f6) : $signed(_GEN_2407); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2409 = 11'h168 == cnt[10:0] ? $signed(-32'sh864c) : $signed(_GEN_2408); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2410 = 11'h169 == cnt[10:0] ? $signed(-32'sh86a1) : $signed(_GEN_2409); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2411 = 11'h16a == cnt[10:0] ? $signed(-32'sh86f7) : $signed(_GEN_2410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2412 = 11'h16b == cnt[10:0] ? $signed(-32'sh874c) : $signed(_GEN_2411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2413 = 11'h16c == cnt[10:0] ? $signed(-32'sh87a1) : $signed(_GEN_2412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2414 = 11'h16d == cnt[10:0] ? $signed(-32'sh87f6) : $signed(_GEN_2413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2415 = 11'h16e == cnt[10:0] ? $signed(-32'sh884c) : $signed(_GEN_2414); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2416 = 11'h16f == cnt[10:0] ? $signed(-32'sh88a1) : $signed(_GEN_2415); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2417 = 11'h170 == cnt[10:0] ? $signed(-32'sh88f6) : $signed(_GEN_2416); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2418 = 11'h171 == cnt[10:0] ? $signed(-32'sh894a) : $signed(_GEN_2417); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2419 = 11'h172 == cnt[10:0] ? $signed(-32'sh899f) : $signed(_GEN_2418); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2420 = 11'h173 == cnt[10:0] ? $signed(-32'sh89f4) : $signed(_GEN_2419); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2421 = 11'h174 == cnt[10:0] ? $signed(-32'sh8a49) : $signed(_GEN_2420); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2422 = 11'h175 == cnt[10:0] ? $signed(-32'sh8a9d) : $signed(_GEN_2421); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2423 = 11'h176 == cnt[10:0] ? $signed(-32'sh8af2) : $signed(_GEN_2422); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2424 = 11'h177 == cnt[10:0] ? $signed(-32'sh8b46) : $signed(_GEN_2423); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2425 = 11'h178 == cnt[10:0] ? $signed(-32'sh8b9a) : $signed(_GEN_2424); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2426 = 11'h179 == cnt[10:0] ? $signed(-32'sh8bef) : $signed(_GEN_2425); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2427 = 11'h17a == cnt[10:0] ? $signed(-32'sh8c43) : $signed(_GEN_2426); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2428 = 11'h17b == cnt[10:0] ? $signed(-32'sh8c97) : $signed(_GEN_2427); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2429 = 11'h17c == cnt[10:0] ? $signed(-32'sh8ceb) : $signed(_GEN_2428); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2430 = 11'h17d == cnt[10:0] ? $signed(-32'sh8d3f) : $signed(_GEN_2429); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2431 = 11'h17e == cnt[10:0] ? $signed(-32'sh8d93) : $signed(_GEN_2430); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2432 = 11'h17f == cnt[10:0] ? $signed(-32'sh8de6) : $signed(_GEN_2431); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2433 = 11'h180 == cnt[10:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2432); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2434 = 11'h181 == cnt[10:0] ? $signed(-32'sh8e8d) : $signed(_GEN_2433); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2435 = 11'h182 == cnt[10:0] ? $signed(-32'sh8ee1) : $signed(_GEN_2434); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2436 = 11'h183 == cnt[10:0] ? $signed(-32'sh8f34) : $signed(_GEN_2435); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2437 = 11'h184 == cnt[10:0] ? $signed(-32'sh8f88) : $signed(_GEN_2436); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2438 = 11'h185 == cnt[10:0] ? $signed(-32'sh8fdb) : $signed(_GEN_2437); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2439 = 11'h186 == cnt[10:0] ? $signed(-32'sh902e) : $signed(_GEN_2438); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2440 = 11'h187 == cnt[10:0] ? $signed(-32'sh9081) : $signed(_GEN_2439); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2441 = 11'h188 == cnt[10:0] ? $signed(-32'sh90d4) : $signed(_GEN_2440); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2442 = 11'h189 == cnt[10:0] ? $signed(-32'sh9127) : $signed(_GEN_2441); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2443 = 11'h18a == cnt[10:0] ? $signed(-32'sh9179) : $signed(_GEN_2442); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2444 = 11'h18b == cnt[10:0] ? $signed(-32'sh91cc) : $signed(_GEN_2443); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2445 = 11'h18c == cnt[10:0] ? $signed(-32'sh921f) : $signed(_GEN_2444); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2446 = 11'h18d == cnt[10:0] ? $signed(-32'sh9271) : $signed(_GEN_2445); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2447 = 11'h18e == cnt[10:0] ? $signed(-32'sh92c4) : $signed(_GEN_2446); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2448 = 11'h18f == cnt[10:0] ? $signed(-32'sh9316) : $signed(_GEN_2447); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2449 = 11'h190 == cnt[10:0] ? $signed(-32'sh9368) : $signed(_GEN_2448); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2450 = 11'h191 == cnt[10:0] ? $signed(-32'sh93ba) : $signed(_GEN_2449); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2451 = 11'h192 == cnt[10:0] ? $signed(-32'sh940c) : $signed(_GEN_2450); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2452 = 11'h193 == cnt[10:0] ? $signed(-32'sh945e) : $signed(_GEN_2451); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2453 = 11'h194 == cnt[10:0] ? $signed(-32'sh94b0) : $signed(_GEN_2452); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2454 = 11'h195 == cnt[10:0] ? $signed(-32'sh9502) : $signed(_GEN_2453); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2455 = 11'h196 == cnt[10:0] ? $signed(-32'sh9554) : $signed(_GEN_2454); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2456 = 11'h197 == cnt[10:0] ? $signed(-32'sh95a5) : $signed(_GEN_2455); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2457 = 11'h198 == cnt[10:0] ? $signed(-32'sh95f7) : $signed(_GEN_2456); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2458 = 11'h199 == cnt[10:0] ? $signed(-32'sh9648) : $signed(_GEN_2457); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2459 = 11'h19a == cnt[10:0] ? $signed(-32'sh969a) : $signed(_GEN_2458); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2460 = 11'h19b == cnt[10:0] ? $signed(-32'sh96eb) : $signed(_GEN_2459); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2461 = 11'h19c == cnt[10:0] ? $signed(-32'sh973c) : $signed(_GEN_2460); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2462 = 11'h19d == cnt[10:0] ? $signed(-32'sh978d) : $signed(_GEN_2461); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2463 = 11'h19e == cnt[10:0] ? $signed(-32'sh97de) : $signed(_GEN_2462); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2464 = 11'h19f == cnt[10:0] ? $signed(-32'sh982f) : $signed(_GEN_2463); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2465 = 11'h1a0 == cnt[10:0] ? $signed(-32'sh9880) : $signed(_GEN_2464); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2466 = 11'h1a1 == cnt[10:0] ? $signed(-32'sh98d0) : $signed(_GEN_2465); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2467 = 11'h1a2 == cnt[10:0] ? $signed(-32'sh9921) : $signed(_GEN_2466); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2468 = 11'h1a3 == cnt[10:0] ? $signed(-32'sh9972) : $signed(_GEN_2467); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2469 = 11'h1a4 == cnt[10:0] ? $signed(-32'sh99c2) : $signed(_GEN_2468); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2470 = 11'h1a5 == cnt[10:0] ? $signed(-32'sh9a12) : $signed(_GEN_2469); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2471 = 11'h1a6 == cnt[10:0] ? $signed(-32'sh9a63) : $signed(_GEN_2470); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2472 = 11'h1a7 == cnt[10:0] ? $signed(-32'sh9ab3) : $signed(_GEN_2471); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2473 = 11'h1a8 == cnt[10:0] ? $signed(-32'sh9b03) : $signed(_GEN_2472); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2474 = 11'h1a9 == cnt[10:0] ? $signed(-32'sh9b53) : $signed(_GEN_2473); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2475 = 11'h1aa == cnt[10:0] ? $signed(-32'sh9ba3) : $signed(_GEN_2474); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2476 = 11'h1ab == cnt[10:0] ? $signed(-32'sh9bf2) : $signed(_GEN_2475); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2477 = 11'h1ac == cnt[10:0] ? $signed(-32'sh9c42) : $signed(_GEN_2476); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2478 = 11'h1ad == cnt[10:0] ? $signed(-32'sh9c92) : $signed(_GEN_2477); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2479 = 11'h1ae == cnt[10:0] ? $signed(-32'sh9ce1) : $signed(_GEN_2478); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2480 = 11'h1af == cnt[10:0] ? $signed(-32'sh9d31) : $signed(_GEN_2479); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2481 = 11'h1b0 == cnt[10:0] ? $signed(-32'sh9d80) : $signed(_GEN_2480); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2482 = 11'h1b1 == cnt[10:0] ? $signed(-32'sh9dcf) : $signed(_GEN_2481); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2483 = 11'h1b2 == cnt[10:0] ? $signed(-32'sh9e1e) : $signed(_GEN_2482); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2484 = 11'h1b3 == cnt[10:0] ? $signed(-32'sh9e6d) : $signed(_GEN_2483); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2485 = 11'h1b4 == cnt[10:0] ? $signed(-32'sh9ebc) : $signed(_GEN_2484); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2486 = 11'h1b5 == cnt[10:0] ? $signed(-32'sh9f0b) : $signed(_GEN_2485); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2487 = 11'h1b6 == cnt[10:0] ? $signed(-32'sh9f5a) : $signed(_GEN_2486); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2488 = 11'h1b7 == cnt[10:0] ? $signed(-32'sh9fa8) : $signed(_GEN_2487); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2489 = 11'h1b8 == cnt[10:0] ? $signed(-32'sh9ff7) : $signed(_GEN_2488); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2490 = 11'h1b9 == cnt[10:0] ? $signed(-32'sha045) : $signed(_GEN_2489); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2491 = 11'h1ba == cnt[10:0] ? $signed(-32'sha094) : $signed(_GEN_2490); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2492 = 11'h1bb == cnt[10:0] ? $signed(-32'sha0e2) : $signed(_GEN_2491); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2493 = 11'h1bc == cnt[10:0] ? $signed(-32'sha130) : $signed(_GEN_2492); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2494 = 11'h1bd == cnt[10:0] ? $signed(-32'sha17e) : $signed(_GEN_2493); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2495 = 11'h1be == cnt[10:0] ? $signed(-32'sha1cc) : $signed(_GEN_2494); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2496 = 11'h1bf == cnt[10:0] ? $signed(-32'sha21a) : $signed(_GEN_2495); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2497 = 11'h1c0 == cnt[10:0] ? $signed(-32'sha268) : $signed(_GEN_2496); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2498 = 11'h1c1 == cnt[10:0] ? $signed(-32'sha2b5) : $signed(_GEN_2497); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2499 = 11'h1c2 == cnt[10:0] ? $signed(-32'sha303) : $signed(_GEN_2498); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2500 = 11'h1c3 == cnt[10:0] ? $signed(-32'sha350) : $signed(_GEN_2499); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2501 = 11'h1c4 == cnt[10:0] ? $signed(-32'sha39e) : $signed(_GEN_2500); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2502 = 11'h1c5 == cnt[10:0] ? $signed(-32'sha3eb) : $signed(_GEN_2501); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2503 = 11'h1c6 == cnt[10:0] ? $signed(-32'sha438) : $signed(_GEN_2502); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2504 = 11'h1c7 == cnt[10:0] ? $signed(-32'sha485) : $signed(_GEN_2503); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2505 = 11'h1c8 == cnt[10:0] ? $signed(-32'sha4d2) : $signed(_GEN_2504); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2506 = 11'h1c9 == cnt[10:0] ? $signed(-32'sha51f) : $signed(_GEN_2505); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2507 = 11'h1ca == cnt[10:0] ? $signed(-32'sha56c) : $signed(_GEN_2506); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2508 = 11'h1cb == cnt[10:0] ? $signed(-32'sha5b8) : $signed(_GEN_2507); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2509 = 11'h1cc == cnt[10:0] ? $signed(-32'sha605) : $signed(_GEN_2508); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2510 = 11'h1cd == cnt[10:0] ? $signed(-32'sha652) : $signed(_GEN_2509); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2511 = 11'h1ce == cnt[10:0] ? $signed(-32'sha69e) : $signed(_GEN_2510); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2512 = 11'h1cf == cnt[10:0] ? $signed(-32'sha6ea) : $signed(_GEN_2511); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2513 = 11'h1d0 == cnt[10:0] ? $signed(-32'sha736) : $signed(_GEN_2512); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2514 = 11'h1d1 == cnt[10:0] ? $signed(-32'sha782) : $signed(_GEN_2513); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2515 = 11'h1d2 == cnt[10:0] ? $signed(-32'sha7ce) : $signed(_GEN_2514); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2516 = 11'h1d3 == cnt[10:0] ? $signed(-32'sha81a) : $signed(_GEN_2515); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2517 = 11'h1d4 == cnt[10:0] ? $signed(-32'sha866) : $signed(_GEN_2516); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2518 = 11'h1d5 == cnt[10:0] ? $signed(-32'sha8b2) : $signed(_GEN_2517); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2519 = 11'h1d6 == cnt[10:0] ? $signed(-32'sha8fd) : $signed(_GEN_2518); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2520 = 11'h1d7 == cnt[10:0] ? $signed(-32'sha949) : $signed(_GEN_2519); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2521 = 11'h1d8 == cnt[10:0] ? $signed(-32'sha994) : $signed(_GEN_2520); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2522 = 11'h1d9 == cnt[10:0] ? $signed(-32'sha9df) : $signed(_GEN_2521); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2523 = 11'h1da == cnt[10:0] ? $signed(-32'shaa2a) : $signed(_GEN_2522); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2524 = 11'h1db == cnt[10:0] ? $signed(-32'shaa76) : $signed(_GEN_2523); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2525 = 11'h1dc == cnt[10:0] ? $signed(-32'shaac1) : $signed(_GEN_2524); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2526 = 11'h1dd == cnt[10:0] ? $signed(-32'shab0b) : $signed(_GEN_2525); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2527 = 11'h1de == cnt[10:0] ? $signed(-32'shab56) : $signed(_GEN_2526); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2528 = 11'h1df == cnt[10:0] ? $signed(-32'shaba1) : $signed(_GEN_2527); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2529 = 11'h1e0 == cnt[10:0] ? $signed(-32'shabeb) : $signed(_GEN_2528); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2530 = 11'h1e1 == cnt[10:0] ? $signed(-32'shac36) : $signed(_GEN_2529); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2531 = 11'h1e2 == cnt[10:0] ? $signed(-32'shac80) : $signed(_GEN_2530); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2532 = 11'h1e3 == cnt[10:0] ? $signed(-32'shacca) : $signed(_GEN_2531); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2533 = 11'h1e4 == cnt[10:0] ? $signed(-32'shad14) : $signed(_GEN_2532); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2534 = 11'h1e5 == cnt[10:0] ? $signed(-32'shad5e) : $signed(_GEN_2533); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2535 = 11'h1e6 == cnt[10:0] ? $signed(-32'shada8) : $signed(_GEN_2534); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2536 = 11'h1e7 == cnt[10:0] ? $signed(-32'shadf2) : $signed(_GEN_2535); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2537 = 11'h1e8 == cnt[10:0] ? $signed(-32'shae3c) : $signed(_GEN_2536); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2538 = 11'h1e9 == cnt[10:0] ? $signed(-32'shae85) : $signed(_GEN_2537); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2539 = 11'h1ea == cnt[10:0] ? $signed(-32'shaecf) : $signed(_GEN_2538); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2540 = 11'h1eb == cnt[10:0] ? $signed(-32'shaf18) : $signed(_GEN_2539); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2541 = 11'h1ec == cnt[10:0] ? $signed(-32'shaf62) : $signed(_GEN_2540); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2542 = 11'h1ed == cnt[10:0] ? $signed(-32'shafab) : $signed(_GEN_2541); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2543 = 11'h1ee == cnt[10:0] ? $signed(-32'shaff4) : $signed(_GEN_2542); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2544 = 11'h1ef == cnt[10:0] ? $signed(-32'shb03d) : $signed(_GEN_2543); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2545 = 11'h1f0 == cnt[10:0] ? $signed(-32'shb086) : $signed(_GEN_2544); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2546 = 11'h1f1 == cnt[10:0] ? $signed(-32'shb0ce) : $signed(_GEN_2545); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2547 = 11'h1f2 == cnt[10:0] ? $signed(-32'shb117) : $signed(_GEN_2546); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2548 = 11'h1f3 == cnt[10:0] ? $signed(-32'shb160) : $signed(_GEN_2547); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2549 = 11'h1f4 == cnt[10:0] ? $signed(-32'shb1a8) : $signed(_GEN_2548); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2550 = 11'h1f5 == cnt[10:0] ? $signed(-32'shb1f0) : $signed(_GEN_2549); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2551 = 11'h1f6 == cnt[10:0] ? $signed(-32'shb239) : $signed(_GEN_2550); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2552 = 11'h1f7 == cnt[10:0] ? $signed(-32'shb281) : $signed(_GEN_2551); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2553 = 11'h1f8 == cnt[10:0] ? $signed(-32'shb2c9) : $signed(_GEN_2552); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2554 = 11'h1f9 == cnt[10:0] ? $signed(-32'shb311) : $signed(_GEN_2553); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2555 = 11'h1fa == cnt[10:0] ? $signed(-32'shb358) : $signed(_GEN_2554); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2556 = 11'h1fb == cnt[10:0] ? $signed(-32'shb3a0) : $signed(_GEN_2555); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2557 = 11'h1fc == cnt[10:0] ? $signed(-32'shb3e8) : $signed(_GEN_2556); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2558 = 11'h1fd == cnt[10:0] ? $signed(-32'shb42f) : $signed(_GEN_2557); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2559 = 11'h1fe == cnt[10:0] ? $signed(-32'shb477) : $signed(_GEN_2558); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2560 = 11'h1ff == cnt[10:0] ? $signed(-32'shb4be) : $signed(_GEN_2559); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2561 = 11'h200 == cnt[10:0] ? $signed(-32'shb505) : $signed(_GEN_2560); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2562 = 11'h201 == cnt[10:0] ? $signed(-32'shb54c) : $signed(_GEN_2561); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2563 = 11'h202 == cnt[10:0] ? $signed(-32'shb593) : $signed(_GEN_2562); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2564 = 11'h203 == cnt[10:0] ? $signed(-32'shb5da) : $signed(_GEN_2563); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2565 = 11'h204 == cnt[10:0] ? $signed(-32'shb620) : $signed(_GEN_2564); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2566 = 11'h205 == cnt[10:0] ? $signed(-32'shb667) : $signed(_GEN_2565); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2567 = 11'h206 == cnt[10:0] ? $signed(-32'shb6ad) : $signed(_GEN_2566); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2568 = 11'h207 == cnt[10:0] ? $signed(-32'shb6f4) : $signed(_GEN_2567); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2569 = 11'h208 == cnt[10:0] ? $signed(-32'shb73a) : $signed(_GEN_2568); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2570 = 11'h209 == cnt[10:0] ? $signed(-32'shb780) : $signed(_GEN_2569); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2571 = 11'h20a == cnt[10:0] ? $signed(-32'shb7c6) : $signed(_GEN_2570); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2572 = 11'h20b == cnt[10:0] ? $signed(-32'shb80c) : $signed(_GEN_2571); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2573 = 11'h20c == cnt[10:0] ? $signed(-32'shb852) : $signed(_GEN_2572); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2574 = 11'h20d == cnt[10:0] ? $signed(-32'shb898) : $signed(_GEN_2573); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2575 = 11'h20e == cnt[10:0] ? $signed(-32'shb8dd) : $signed(_GEN_2574); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2576 = 11'h20f == cnt[10:0] ? $signed(-32'shb923) : $signed(_GEN_2575); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2577 = 11'h210 == cnt[10:0] ? $signed(-32'shb968) : $signed(_GEN_2576); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2578 = 11'h211 == cnt[10:0] ? $signed(-32'shb9ae) : $signed(_GEN_2577); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2579 = 11'h212 == cnt[10:0] ? $signed(-32'shb9f3) : $signed(_GEN_2578); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2580 = 11'h213 == cnt[10:0] ? $signed(-32'shba38) : $signed(_GEN_2579); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2581 = 11'h214 == cnt[10:0] ? $signed(-32'shba7d) : $signed(_GEN_2580); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2582 = 11'h215 == cnt[10:0] ? $signed(-32'shbac1) : $signed(_GEN_2581); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2583 = 11'h216 == cnt[10:0] ? $signed(-32'shbb06) : $signed(_GEN_2582); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2584 = 11'h217 == cnt[10:0] ? $signed(-32'shbb4b) : $signed(_GEN_2583); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2585 = 11'h218 == cnt[10:0] ? $signed(-32'shbb8f) : $signed(_GEN_2584); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2586 = 11'h219 == cnt[10:0] ? $signed(-32'shbbd4) : $signed(_GEN_2585); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2587 = 11'h21a == cnt[10:0] ? $signed(-32'shbc18) : $signed(_GEN_2586); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2588 = 11'h21b == cnt[10:0] ? $signed(-32'shbc5c) : $signed(_GEN_2587); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2589 = 11'h21c == cnt[10:0] ? $signed(-32'shbca0) : $signed(_GEN_2588); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2590 = 11'h21d == cnt[10:0] ? $signed(-32'shbce4) : $signed(_GEN_2589); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2591 = 11'h21e == cnt[10:0] ? $signed(-32'shbd28) : $signed(_GEN_2590); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2592 = 11'h21f == cnt[10:0] ? $signed(-32'shbd6b) : $signed(_GEN_2591); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2593 = 11'h220 == cnt[10:0] ? $signed(-32'shbdaf) : $signed(_GEN_2592); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2594 = 11'h221 == cnt[10:0] ? $signed(-32'shbdf2) : $signed(_GEN_2593); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2595 = 11'h222 == cnt[10:0] ? $signed(-32'shbe36) : $signed(_GEN_2594); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2596 = 11'h223 == cnt[10:0] ? $signed(-32'shbe79) : $signed(_GEN_2595); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2597 = 11'h224 == cnt[10:0] ? $signed(-32'shbebc) : $signed(_GEN_2596); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2598 = 11'h225 == cnt[10:0] ? $signed(-32'shbeff) : $signed(_GEN_2597); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2599 = 11'h226 == cnt[10:0] ? $signed(-32'shbf42) : $signed(_GEN_2598); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2600 = 11'h227 == cnt[10:0] ? $signed(-32'shbf85) : $signed(_GEN_2599); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2601 = 11'h228 == cnt[10:0] ? $signed(-32'shbfc7) : $signed(_GEN_2600); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2602 = 11'h229 == cnt[10:0] ? $signed(-32'shc00a) : $signed(_GEN_2601); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2603 = 11'h22a == cnt[10:0] ? $signed(-32'shc04c) : $signed(_GEN_2602); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2604 = 11'h22b == cnt[10:0] ? $signed(-32'shc08f) : $signed(_GEN_2603); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2605 = 11'h22c == cnt[10:0] ? $signed(-32'shc0d1) : $signed(_GEN_2604); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2606 = 11'h22d == cnt[10:0] ? $signed(-32'shc113) : $signed(_GEN_2605); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2607 = 11'h22e == cnt[10:0] ? $signed(-32'shc155) : $signed(_GEN_2606); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2608 = 11'h22f == cnt[10:0] ? $signed(-32'shc197) : $signed(_GEN_2607); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2609 = 11'h230 == cnt[10:0] ? $signed(-32'shc1d8) : $signed(_GEN_2608); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2610 = 11'h231 == cnt[10:0] ? $signed(-32'shc21a) : $signed(_GEN_2609); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2611 = 11'h232 == cnt[10:0] ? $signed(-32'shc25c) : $signed(_GEN_2610); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2612 = 11'h233 == cnt[10:0] ? $signed(-32'shc29d) : $signed(_GEN_2611); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2613 = 11'h234 == cnt[10:0] ? $signed(-32'shc2de) : $signed(_GEN_2612); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2614 = 11'h235 == cnt[10:0] ? $signed(-32'shc31f) : $signed(_GEN_2613); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2615 = 11'h236 == cnt[10:0] ? $signed(-32'shc360) : $signed(_GEN_2614); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2616 = 11'h237 == cnt[10:0] ? $signed(-32'shc3a1) : $signed(_GEN_2615); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2617 = 11'h238 == cnt[10:0] ? $signed(-32'shc3e2) : $signed(_GEN_2616); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2618 = 11'h239 == cnt[10:0] ? $signed(-32'shc423) : $signed(_GEN_2617); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2619 = 11'h23a == cnt[10:0] ? $signed(-32'shc463) : $signed(_GEN_2618); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2620 = 11'h23b == cnt[10:0] ? $signed(-32'shc4a4) : $signed(_GEN_2619); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2621 = 11'h23c == cnt[10:0] ? $signed(-32'shc4e4) : $signed(_GEN_2620); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2622 = 11'h23d == cnt[10:0] ? $signed(-32'shc524) : $signed(_GEN_2621); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2623 = 11'h23e == cnt[10:0] ? $signed(-32'shc564) : $signed(_GEN_2622); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2624 = 11'h23f == cnt[10:0] ? $signed(-32'shc5a4) : $signed(_GEN_2623); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2625 = 11'h240 == cnt[10:0] ? $signed(-32'shc5e4) : $signed(_GEN_2624); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2626 = 11'h241 == cnt[10:0] ? $signed(-32'shc624) : $signed(_GEN_2625); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2627 = 11'h242 == cnt[10:0] ? $signed(-32'shc663) : $signed(_GEN_2626); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2628 = 11'h243 == cnt[10:0] ? $signed(-32'shc6a3) : $signed(_GEN_2627); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2629 = 11'h244 == cnt[10:0] ? $signed(-32'shc6e2) : $signed(_GEN_2628); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2630 = 11'h245 == cnt[10:0] ? $signed(-32'shc721) : $signed(_GEN_2629); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2631 = 11'h246 == cnt[10:0] ? $signed(-32'shc761) : $signed(_GEN_2630); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2632 = 11'h247 == cnt[10:0] ? $signed(-32'shc7a0) : $signed(_GEN_2631); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2633 = 11'h248 == cnt[10:0] ? $signed(-32'shc7de) : $signed(_GEN_2632); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2634 = 11'h249 == cnt[10:0] ? $signed(-32'shc81d) : $signed(_GEN_2633); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2635 = 11'h24a == cnt[10:0] ? $signed(-32'shc85c) : $signed(_GEN_2634); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2636 = 11'h24b == cnt[10:0] ? $signed(-32'shc89a) : $signed(_GEN_2635); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2637 = 11'h24c == cnt[10:0] ? $signed(-32'shc8d9) : $signed(_GEN_2636); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2638 = 11'h24d == cnt[10:0] ? $signed(-32'shc917) : $signed(_GEN_2637); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2639 = 11'h24e == cnt[10:0] ? $signed(-32'shc955) : $signed(_GEN_2638); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2640 = 11'h24f == cnt[10:0] ? $signed(-32'shc993) : $signed(_GEN_2639); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2641 = 11'h250 == cnt[10:0] ? $signed(-32'shc9d1) : $signed(_GEN_2640); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2642 = 11'h251 == cnt[10:0] ? $signed(-32'shca0f) : $signed(_GEN_2641); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2643 = 11'h252 == cnt[10:0] ? $signed(-32'shca4d) : $signed(_GEN_2642); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2644 = 11'h253 == cnt[10:0] ? $signed(-32'shca8a) : $signed(_GEN_2643); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2645 = 11'h254 == cnt[10:0] ? $signed(-32'shcac7) : $signed(_GEN_2644); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2646 = 11'h255 == cnt[10:0] ? $signed(-32'shcb05) : $signed(_GEN_2645); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2647 = 11'h256 == cnt[10:0] ? $signed(-32'shcb42) : $signed(_GEN_2646); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2648 = 11'h257 == cnt[10:0] ? $signed(-32'shcb7f) : $signed(_GEN_2647); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2649 = 11'h258 == cnt[10:0] ? $signed(-32'shcbbc) : $signed(_GEN_2648); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2650 = 11'h259 == cnt[10:0] ? $signed(-32'shcbf9) : $signed(_GEN_2649); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2651 = 11'h25a == cnt[10:0] ? $signed(-32'shcc35) : $signed(_GEN_2650); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2652 = 11'h25b == cnt[10:0] ? $signed(-32'shcc72) : $signed(_GEN_2651); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2653 = 11'h25c == cnt[10:0] ? $signed(-32'shccae) : $signed(_GEN_2652); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2654 = 11'h25d == cnt[10:0] ? $signed(-32'shcceb) : $signed(_GEN_2653); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2655 = 11'h25e == cnt[10:0] ? $signed(-32'shcd27) : $signed(_GEN_2654); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2656 = 11'h25f == cnt[10:0] ? $signed(-32'shcd63) : $signed(_GEN_2655); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2657 = 11'h260 == cnt[10:0] ? $signed(-32'shcd9f) : $signed(_GEN_2656); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2658 = 11'h261 == cnt[10:0] ? $signed(-32'shcddb) : $signed(_GEN_2657); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2659 = 11'h262 == cnt[10:0] ? $signed(-32'shce17) : $signed(_GEN_2658); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2660 = 11'h263 == cnt[10:0] ? $signed(-32'shce52) : $signed(_GEN_2659); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2661 = 11'h264 == cnt[10:0] ? $signed(-32'shce8e) : $signed(_GEN_2660); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2662 = 11'h265 == cnt[10:0] ? $signed(-32'shcec9) : $signed(_GEN_2661); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2663 = 11'h266 == cnt[10:0] ? $signed(-32'shcf04) : $signed(_GEN_2662); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2664 = 11'h267 == cnt[10:0] ? $signed(-32'shcf3f) : $signed(_GEN_2663); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2665 = 11'h268 == cnt[10:0] ? $signed(-32'shcf7a) : $signed(_GEN_2664); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2666 = 11'h269 == cnt[10:0] ? $signed(-32'shcfb5) : $signed(_GEN_2665); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2667 = 11'h26a == cnt[10:0] ? $signed(-32'shcff0) : $signed(_GEN_2666); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2668 = 11'h26b == cnt[10:0] ? $signed(-32'shd02a) : $signed(_GEN_2667); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2669 = 11'h26c == cnt[10:0] ? $signed(-32'shd065) : $signed(_GEN_2668); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2670 = 11'h26d == cnt[10:0] ? $signed(-32'shd09f) : $signed(_GEN_2669); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2671 = 11'h26e == cnt[10:0] ? $signed(-32'shd0d9) : $signed(_GEN_2670); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2672 = 11'h26f == cnt[10:0] ? $signed(-32'shd113) : $signed(_GEN_2671); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2673 = 11'h270 == cnt[10:0] ? $signed(-32'shd14d) : $signed(_GEN_2672); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2674 = 11'h271 == cnt[10:0] ? $signed(-32'shd187) : $signed(_GEN_2673); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2675 = 11'h272 == cnt[10:0] ? $signed(-32'shd1c1) : $signed(_GEN_2674); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2676 = 11'h273 == cnt[10:0] ? $signed(-32'shd1fa) : $signed(_GEN_2675); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2677 = 11'h274 == cnt[10:0] ? $signed(-32'shd234) : $signed(_GEN_2676); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2678 = 11'h275 == cnt[10:0] ? $signed(-32'shd26d) : $signed(_GEN_2677); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2679 = 11'h276 == cnt[10:0] ? $signed(-32'shd2a6) : $signed(_GEN_2678); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2680 = 11'h277 == cnt[10:0] ? $signed(-32'shd2df) : $signed(_GEN_2679); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2681 = 11'h278 == cnt[10:0] ? $signed(-32'shd318) : $signed(_GEN_2680); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2682 = 11'h279 == cnt[10:0] ? $signed(-32'shd351) : $signed(_GEN_2681); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2683 = 11'h27a == cnt[10:0] ? $signed(-32'shd38a) : $signed(_GEN_2682); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2684 = 11'h27b == cnt[10:0] ? $signed(-32'shd3c2) : $signed(_GEN_2683); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2685 = 11'h27c == cnt[10:0] ? $signed(-32'shd3fb) : $signed(_GEN_2684); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2686 = 11'h27d == cnt[10:0] ? $signed(-32'shd433) : $signed(_GEN_2685); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2687 = 11'h27e == cnt[10:0] ? $signed(-32'shd46b) : $signed(_GEN_2686); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2688 = 11'h27f == cnt[10:0] ? $signed(-32'shd4a3) : $signed(_GEN_2687); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2689 = 11'h280 == cnt[10:0] ? $signed(-32'shd4db) : $signed(_GEN_2688); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2690 = 11'h281 == cnt[10:0] ? $signed(-32'shd513) : $signed(_GEN_2689); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2691 = 11'h282 == cnt[10:0] ? $signed(-32'shd54b) : $signed(_GEN_2690); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2692 = 11'h283 == cnt[10:0] ? $signed(-32'shd582) : $signed(_GEN_2691); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2693 = 11'h284 == cnt[10:0] ? $signed(-32'shd5ba) : $signed(_GEN_2692); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2694 = 11'h285 == cnt[10:0] ? $signed(-32'shd5f1) : $signed(_GEN_2693); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2695 = 11'h286 == cnt[10:0] ? $signed(-32'shd628) : $signed(_GEN_2694); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2696 = 11'h287 == cnt[10:0] ? $signed(-32'shd65f) : $signed(_GEN_2695); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2697 = 11'h288 == cnt[10:0] ? $signed(-32'shd696) : $signed(_GEN_2696); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2698 = 11'h289 == cnt[10:0] ? $signed(-32'shd6cd) : $signed(_GEN_2697); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2699 = 11'h28a == cnt[10:0] ? $signed(-32'shd703) : $signed(_GEN_2698); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2700 = 11'h28b == cnt[10:0] ? $signed(-32'shd73a) : $signed(_GEN_2699); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2701 = 11'h28c == cnt[10:0] ? $signed(-32'shd770) : $signed(_GEN_2700); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2702 = 11'h28d == cnt[10:0] ? $signed(-32'shd7a6) : $signed(_GEN_2701); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2703 = 11'h28e == cnt[10:0] ? $signed(-32'shd7dc) : $signed(_GEN_2702); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2704 = 11'h28f == cnt[10:0] ? $signed(-32'shd812) : $signed(_GEN_2703); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2705 = 11'h290 == cnt[10:0] ? $signed(-32'shd848) : $signed(_GEN_2704); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2706 = 11'h291 == cnt[10:0] ? $signed(-32'shd87e) : $signed(_GEN_2705); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2707 = 11'h292 == cnt[10:0] ? $signed(-32'shd8b4) : $signed(_GEN_2706); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2708 = 11'h293 == cnt[10:0] ? $signed(-32'shd8e9) : $signed(_GEN_2707); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2709 = 11'h294 == cnt[10:0] ? $signed(-32'shd91e) : $signed(_GEN_2708); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2710 = 11'h295 == cnt[10:0] ? $signed(-32'shd954) : $signed(_GEN_2709); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2711 = 11'h296 == cnt[10:0] ? $signed(-32'shd989) : $signed(_GEN_2710); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2712 = 11'h297 == cnt[10:0] ? $signed(-32'shd9be) : $signed(_GEN_2711); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2713 = 11'h298 == cnt[10:0] ? $signed(-32'shd9f2) : $signed(_GEN_2712); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2714 = 11'h299 == cnt[10:0] ? $signed(-32'shda27) : $signed(_GEN_2713); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2715 = 11'h29a == cnt[10:0] ? $signed(-32'shda5c) : $signed(_GEN_2714); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2716 = 11'h29b == cnt[10:0] ? $signed(-32'shda90) : $signed(_GEN_2715); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2717 = 11'h29c == cnt[10:0] ? $signed(-32'shdac4) : $signed(_GEN_2716); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2718 = 11'h29d == cnt[10:0] ? $signed(-32'shdaf8) : $signed(_GEN_2717); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2719 = 11'h29e == cnt[10:0] ? $signed(-32'shdb2c) : $signed(_GEN_2718); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2720 = 11'h29f == cnt[10:0] ? $signed(-32'shdb60) : $signed(_GEN_2719); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2721 = 11'h2a0 == cnt[10:0] ? $signed(-32'shdb94) : $signed(_GEN_2720); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2722 = 11'h2a1 == cnt[10:0] ? $signed(-32'shdbc8) : $signed(_GEN_2721); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2723 = 11'h2a2 == cnt[10:0] ? $signed(-32'shdbfb) : $signed(_GEN_2722); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2724 = 11'h2a3 == cnt[10:0] ? $signed(-32'shdc2f) : $signed(_GEN_2723); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2725 = 11'h2a4 == cnt[10:0] ? $signed(-32'shdc62) : $signed(_GEN_2724); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2726 = 11'h2a5 == cnt[10:0] ? $signed(-32'shdc95) : $signed(_GEN_2725); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2727 = 11'h2a6 == cnt[10:0] ? $signed(-32'shdcc8) : $signed(_GEN_2726); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2728 = 11'h2a7 == cnt[10:0] ? $signed(-32'shdcfb) : $signed(_GEN_2727); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2729 = 11'h2a8 == cnt[10:0] ? $signed(-32'shdd2d) : $signed(_GEN_2728); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2730 = 11'h2a9 == cnt[10:0] ? $signed(-32'shdd60) : $signed(_GEN_2729); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2731 = 11'h2aa == cnt[10:0] ? $signed(-32'shdd92) : $signed(_GEN_2730); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2732 = 11'h2ab == cnt[10:0] ? $signed(-32'shddc5) : $signed(_GEN_2731); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2733 = 11'h2ac == cnt[10:0] ? $signed(-32'shddf7) : $signed(_GEN_2732); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2734 = 11'h2ad == cnt[10:0] ? $signed(-32'shde29) : $signed(_GEN_2733); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2735 = 11'h2ae == cnt[10:0] ? $signed(-32'shde5b) : $signed(_GEN_2734); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2736 = 11'h2af == cnt[10:0] ? $signed(-32'shde8c) : $signed(_GEN_2735); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2737 = 11'h2b0 == cnt[10:0] ? $signed(-32'shdebe) : $signed(_GEN_2736); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2738 = 11'h2b1 == cnt[10:0] ? $signed(-32'shdef0) : $signed(_GEN_2737); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2739 = 11'h2b2 == cnt[10:0] ? $signed(-32'shdf21) : $signed(_GEN_2738); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2740 = 11'h2b3 == cnt[10:0] ? $signed(-32'shdf52) : $signed(_GEN_2739); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2741 = 11'h2b4 == cnt[10:0] ? $signed(-32'shdf83) : $signed(_GEN_2740); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2742 = 11'h2b5 == cnt[10:0] ? $signed(-32'shdfb4) : $signed(_GEN_2741); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2743 = 11'h2b6 == cnt[10:0] ? $signed(-32'shdfe5) : $signed(_GEN_2742); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2744 = 11'h2b7 == cnt[10:0] ? $signed(-32'she016) : $signed(_GEN_2743); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2745 = 11'h2b8 == cnt[10:0] ? $signed(-32'she046) : $signed(_GEN_2744); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2746 = 11'h2b9 == cnt[10:0] ? $signed(-32'she077) : $signed(_GEN_2745); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2747 = 11'h2ba == cnt[10:0] ? $signed(-32'she0a7) : $signed(_GEN_2746); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2748 = 11'h2bb == cnt[10:0] ? $signed(-32'she0d7) : $signed(_GEN_2747); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2749 = 11'h2bc == cnt[10:0] ? $signed(-32'she107) : $signed(_GEN_2748); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2750 = 11'h2bd == cnt[10:0] ? $signed(-32'she137) : $signed(_GEN_2749); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2751 = 11'h2be == cnt[10:0] ? $signed(-32'she167) : $signed(_GEN_2750); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2752 = 11'h2bf == cnt[10:0] ? $signed(-32'she196) : $signed(_GEN_2751); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2753 = 11'h2c0 == cnt[10:0] ? $signed(-32'she1c6) : $signed(_GEN_2752); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2754 = 11'h2c1 == cnt[10:0] ? $signed(-32'she1f5) : $signed(_GEN_2753); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2755 = 11'h2c2 == cnt[10:0] ? $signed(-32'she224) : $signed(_GEN_2754); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2756 = 11'h2c3 == cnt[10:0] ? $signed(-32'she253) : $signed(_GEN_2755); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2757 = 11'h2c4 == cnt[10:0] ? $signed(-32'she282) : $signed(_GEN_2756); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2758 = 11'h2c5 == cnt[10:0] ? $signed(-32'she2b1) : $signed(_GEN_2757); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2759 = 11'h2c6 == cnt[10:0] ? $signed(-32'she2df) : $signed(_GEN_2758); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2760 = 11'h2c7 == cnt[10:0] ? $signed(-32'she30e) : $signed(_GEN_2759); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2761 = 11'h2c8 == cnt[10:0] ? $signed(-32'she33c) : $signed(_GEN_2760); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2762 = 11'h2c9 == cnt[10:0] ? $signed(-32'she36b) : $signed(_GEN_2761); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2763 = 11'h2ca == cnt[10:0] ? $signed(-32'she399) : $signed(_GEN_2762); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2764 = 11'h2cb == cnt[10:0] ? $signed(-32'she3c7) : $signed(_GEN_2763); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2765 = 11'h2cc == cnt[10:0] ? $signed(-32'she3f4) : $signed(_GEN_2764); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2766 = 11'h2cd == cnt[10:0] ? $signed(-32'she422) : $signed(_GEN_2765); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2767 = 11'h2ce == cnt[10:0] ? $signed(-32'she450) : $signed(_GEN_2766); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2768 = 11'h2cf == cnt[10:0] ? $signed(-32'she47d) : $signed(_GEN_2767); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2769 = 11'h2d0 == cnt[10:0] ? $signed(-32'she4aa) : $signed(_GEN_2768); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2770 = 11'h2d1 == cnt[10:0] ? $signed(-32'she4d7) : $signed(_GEN_2769); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2771 = 11'h2d2 == cnt[10:0] ? $signed(-32'she504) : $signed(_GEN_2770); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2772 = 11'h2d3 == cnt[10:0] ? $signed(-32'she531) : $signed(_GEN_2771); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2773 = 11'h2d4 == cnt[10:0] ? $signed(-32'she55e) : $signed(_GEN_2772); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2774 = 11'h2d5 == cnt[10:0] ? $signed(-32'she58b) : $signed(_GEN_2773); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2775 = 11'h2d6 == cnt[10:0] ? $signed(-32'she5b7) : $signed(_GEN_2774); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2776 = 11'h2d7 == cnt[10:0] ? $signed(-32'she5e3) : $signed(_GEN_2775); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2777 = 11'h2d8 == cnt[10:0] ? $signed(-32'she610) : $signed(_GEN_2776); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2778 = 11'h2d9 == cnt[10:0] ? $signed(-32'she63c) : $signed(_GEN_2777); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2779 = 11'h2da == cnt[10:0] ? $signed(-32'she667) : $signed(_GEN_2778); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2780 = 11'h2db == cnt[10:0] ? $signed(-32'she693) : $signed(_GEN_2779); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2781 = 11'h2dc == cnt[10:0] ? $signed(-32'she6bf) : $signed(_GEN_2780); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2782 = 11'h2dd == cnt[10:0] ? $signed(-32'she6ea) : $signed(_GEN_2781); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2783 = 11'h2de == cnt[10:0] ? $signed(-32'she716) : $signed(_GEN_2782); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2784 = 11'h2df == cnt[10:0] ? $signed(-32'she741) : $signed(_GEN_2783); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2785 = 11'h2e0 == cnt[10:0] ? $signed(-32'she76c) : $signed(_GEN_2784); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2786 = 11'h2e1 == cnt[10:0] ? $signed(-32'she797) : $signed(_GEN_2785); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2787 = 11'h2e2 == cnt[10:0] ? $signed(-32'she7c2) : $signed(_GEN_2786); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2788 = 11'h2e3 == cnt[10:0] ? $signed(-32'she7ec) : $signed(_GEN_2787); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2789 = 11'h2e4 == cnt[10:0] ? $signed(-32'she817) : $signed(_GEN_2788); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2790 = 11'h2e5 == cnt[10:0] ? $signed(-32'she841) : $signed(_GEN_2789); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2791 = 11'h2e6 == cnt[10:0] ? $signed(-32'she86b) : $signed(_GEN_2790); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2792 = 11'h2e7 == cnt[10:0] ? $signed(-32'she895) : $signed(_GEN_2791); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2793 = 11'h2e8 == cnt[10:0] ? $signed(-32'she8bf) : $signed(_GEN_2792); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2794 = 11'h2e9 == cnt[10:0] ? $signed(-32'she8e9) : $signed(_GEN_2793); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2795 = 11'h2ea == cnt[10:0] ? $signed(-32'she913) : $signed(_GEN_2794); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2796 = 11'h2eb == cnt[10:0] ? $signed(-32'she93c) : $signed(_GEN_2795); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2797 = 11'h2ec == cnt[10:0] ? $signed(-32'she966) : $signed(_GEN_2796); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2798 = 11'h2ed == cnt[10:0] ? $signed(-32'she98f) : $signed(_GEN_2797); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2799 = 11'h2ee == cnt[10:0] ? $signed(-32'she9b8) : $signed(_GEN_2798); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2800 = 11'h2ef == cnt[10:0] ? $signed(-32'she9e1) : $signed(_GEN_2799); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2801 = 11'h2f0 == cnt[10:0] ? $signed(-32'shea0a) : $signed(_GEN_2800); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2802 = 11'h2f1 == cnt[10:0] ? $signed(-32'shea32) : $signed(_GEN_2801); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2803 = 11'h2f2 == cnt[10:0] ? $signed(-32'shea5b) : $signed(_GEN_2802); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2804 = 11'h2f3 == cnt[10:0] ? $signed(-32'shea83) : $signed(_GEN_2803); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2805 = 11'h2f4 == cnt[10:0] ? $signed(-32'sheaab) : $signed(_GEN_2804); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2806 = 11'h2f5 == cnt[10:0] ? $signed(-32'shead4) : $signed(_GEN_2805); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2807 = 11'h2f6 == cnt[10:0] ? $signed(-32'sheafc) : $signed(_GEN_2806); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2808 = 11'h2f7 == cnt[10:0] ? $signed(-32'sheb23) : $signed(_GEN_2807); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2809 = 11'h2f8 == cnt[10:0] ? $signed(-32'sheb4b) : $signed(_GEN_2808); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2810 = 11'h2f9 == cnt[10:0] ? $signed(-32'sheb73) : $signed(_GEN_2809); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2811 = 11'h2fa == cnt[10:0] ? $signed(-32'sheb9a) : $signed(_GEN_2810); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2812 = 11'h2fb == cnt[10:0] ? $signed(-32'shebc1) : $signed(_GEN_2811); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2813 = 11'h2fc == cnt[10:0] ? $signed(-32'shebe8) : $signed(_GEN_2812); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2814 = 11'h2fd == cnt[10:0] ? $signed(-32'shec0f) : $signed(_GEN_2813); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2815 = 11'h2fe == cnt[10:0] ? $signed(-32'shec36) : $signed(_GEN_2814); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2816 = 11'h2ff == cnt[10:0] ? $signed(-32'shec5d) : $signed(_GEN_2815); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2817 = 11'h300 == cnt[10:0] ? $signed(-32'shec83) : $signed(_GEN_2816); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2818 = 11'h301 == cnt[10:0] ? $signed(-32'shecaa) : $signed(_GEN_2817); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2819 = 11'h302 == cnt[10:0] ? $signed(-32'shecd0) : $signed(_GEN_2818); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2820 = 11'h303 == cnt[10:0] ? $signed(-32'shecf6) : $signed(_GEN_2819); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2821 = 11'h304 == cnt[10:0] ? $signed(-32'shed1c) : $signed(_GEN_2820); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2822 = 11'h305 == cnt[10:0] ? $signed(-32'shed42) : $signed(_GEN_2821); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2823 = 11'h306 == cnt[10:0] ? $signed(-32'shed68) : $signed(_GEN_2822); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2824 = 11'h307 == cnt[10:0] ? $signed(-32'shed8d) : $signed(_GEN_2823); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2825 = 11'h308 == cnt[10:0] ? $signed(-32'shedb3) : $signed(_GEN_2824); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2826 = 11'h309 == cnt[10:0] ? $signed(-32'shedd8) : $signed(_GEN_2825); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2827 = 11'h30a == cnt[10:0] ? $signed(-32'shedfd) : $signed(_GEN_2826); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2828 = 11'h30b == cnt[10:0] ? $signed(-32'shee22) : $signed(_GEN_2827); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2829 = 11'h30c == cnt[10:0] ? $signed(-32'shee47) : $signed(_GEN_2828); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2830 = 11'h30d == cnt[10:0] ? $signed(-32'shee6b) : $signed(_GEN_2829); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2831 = 11'h30e == cnt[10:0] ? $signed(-32'shee90) : $signed(_GEN_2830); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2832 = 11'h30f == cnt[10:0] ? $signed(-32'sheeb4) : $signed(_GEN_2831); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2833 = 11'h310 == cnt[10:0] ? $signed(-32'sheed9) : $signed(_GEN_2832); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2834 = 11'h311 == cnt[10:0] ? $signed(-32'sheefd) : $signed(_GEN_2833); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2835 = 11'h312 == cnt[10:0] ? $signed(-32'shef21) : $signed(_GEN_2834); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2836 = 11'h313 == cnt[10:0] ? $signed(-32'shef45) : $signed(_GEN_2835); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2837 = 11'h314 == cnt[10:0] ? $signed(-32'shef68) : $signed(_GEN_2836); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2838 = 11'h315 == cnt[10:0] ? $signed(-32'shef8c) : $signed(_GEN_2837); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2839 = 11'h316 == cnt[10:0] ? $signed(-32'shefaf) : $signed(_GEN_2838); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2840 = 11'h317 == cnt[10:0] ? $signed(-32'shefd2) : $signed(_GEN_2839); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2841 = 11'h318 == cnt[10:0] ? $signed(-32'sheff5) : $signed(_GEN_2840); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2842 = 11'h319 == cnt[10:0] ? $signed(-32'shf018) : $signed(_GEN_2841); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2843 = 11'h31a == cnt[10:0] ? $signed(-32'shf03b) : $signed(_GEN_2842); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2844 = 11'h31b == cnt[10:0] ? $signed(-32'shf05e) : $signed(_GEN_2843); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2845 = 11'h31c == cnt[10:0] ? $signed(-32'shf080) : $signed(_GEN_2844); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2846 = 11'h31d == cnt[10:0] ? $signed(-32'shf0a3) : $signed(_GEN_2845); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2847 = 11'h31e == cnt[10:0] ? $signed(-32'shf0c5) : $signed(_GEN_2846); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2848 = 11'h31f == cnt[10:0] ? $signed(-32'shf0e7) : $signed(_GEN_2847); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2849 = 11'h320 == cnt[10:0] ? $signed(-32'shf109) : $signed(_GEN_2848); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2850 = 11'h321 == cnt[10:0] ? $signed(-32'shf12b) : $signed(_GEN_2849); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2851 = 11'h322 == cnt[10:0] ? $signed(-32'shf14c) : $signed(_GEN_2850); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2852 = 11'h323 == cnt[10:0] ? $signed(-32'shf16e) : $signed(_GEN_2851); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2853 = 11'h324 == cnt[10:0] ? $signed(-32'shf18f) : $signed(_GEN_2852); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2854 = 11'h325 == cnt[10:0] ? $signed(-32'shf1b1) : $signed(_GEN_2853); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2855 = 11'h326 == cnt[10:0] ? $signed(-32'shf1d2) : $signed(_GEN_2854); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2856 = 11'h327 == cnt[10:0] ? $signed(-32'shf1f3) : $signed(_GEN_2855); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2857 = 11'h328 == cnt[10:0] ? $signed(-32'shf213) : $signed(_GEN_2856); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2858 = 11'h329 == cnt[10:0] ? $signed(-32'shf234) : $signed(_GEN_2857); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2859 = 11'h32a == cnt[10:0] ? $signed(-32'shf254) : $signed(_GEN_2858); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2860 = 11'h32b == cnt[10:0] ? $signed(-32'shf275) : $signed(_GEN_2859); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2861 = 11'h32c == cnt[10:0] ? $signed(-32'shf295) : $signed(_GEN_2860); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2862 = 11'h32d == cnt[10:0] ? $signed(-32'shf2b5) : $signed(_GEN_2861); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2863 = 11'h32e == cnt[10:0] ? $signed(-32'shf2d5) : $signed(_GEN_2862); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2864 = 11'h32f == cnt[10:0] ? $signed(-32'shf2f5) : $signed(_GEN_2863); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2865 = 11'h330 == cnt[10:0] ? $signed(-32'shf314) : $signed(_GEN_2864); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2866 = 11'h331 == cnt[10:0] ? $signed(-32'shf334) : $signed(_GEN_2865); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2867 = 11'h332 == cnt[10:0] ? $signed(-32'shf353) : $signed(_GEN_2866); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2868 = 11'h333 == cnt[10:0] ? $signed(-32'shf372) : $signed(_GEN_2867); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2869 = 11'h334 == cnt[10:0] ? $signed(-32'shf391) : $signed(_GEN_2868); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2870 = 11'h335 == cnt[10:0] ? $signed(-32'shf3b0) : $signed(_GEN_2869); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2871 = 11'h336 == cnt[10:0] ? $signed(-32'shf3cf) : $signed(_GEN_2870); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2872 = 11'h337 == cnt[10:0] ? $signed(-32'shf3ed) : $signed(_GEN_2871); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2873 = 11'h338 == cnt[10:0] ? $signed(-32'shf40c) : $signed(_GEN_2872); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2874 = 11'h339 == cnt[10:0] ? $signed(-32'shf42a) : $signed(_GEN_2873); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2875 = 11'h33a == cnt[10:0] ? $signed(-32'shf448) : $signed(_GEN_2874); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2876 = 11'h33b == cnt[10:0] ? $signed(-32'shf466) : $signed(_GEN_2875); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2877 = 11'h33c == cnt[10:0] ? $signed(-32'shf484) : $signed(_GEN_2876); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2878 = 11'h33d == cnt[10:0] ? $signed(-32'shf4a2) : $signed(_GEN_2877); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2879 = 11'h33e == cnt[10:0] ? $signed(-32'shf4bf) : $signed(_GEN_2878); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2880 = 11'h33f == cnt[10:0] ? $signed(-32'shf4dd) : $signed(_GEN_2879); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2881 = 11'h340 == cnt[10:0] ? $signed(-32'shf4fa) : $signed(_GEN_2880); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2882 = 11'h341 == cnt[10:0] ? $signed(-32'shf517) : $signed(_GEN_2881); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2883 = 11'h342 == cnt[10:0] ? $signed(-32'shf534) : $signed(_GEN_2882); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2884 = 11'h343 == cnt[10:0] ? $signed(-32'shf551) : $signed(_GEN_2883); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2885 = 11'h344 == cnt[10:0] ? $signed(-32'shf56e) : $signed(_GEN_2884); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2886 = 11'h345 == cnt[10:0] ? $signed(-32'shf58a) : $signed(_GEN_2885); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2887 = 11'h346 == cnt[10:0] ? $signed(-32'shf5a6) : $signed(_GEN_2886); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2888 = 11'h347 == cnt[10:0] ? $signed(-32'shf5c3) : $signed(_GEN_2887); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2889 = 11'h348 == cnt[10:0] ? $signed(-32'shf5df) : $signed(_GEN_2888); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2890 = 11'h349 == cnt[10:0] ? $signed(-32'shf5fb) : $signed(_GEN_2889); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2891 = 11'h34a == cnt[10:0] ? $signed(-32'shf616) : $signed(_GEN_2890); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2892 = 11'h34b == cnt[10:0] ? $signed(-32'shf632) : $signed(_GEN_2891); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2893 = 11'h34c == cnt[10:0] ? $signed(-32'shf64e) : $signed(_GEN_2892); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2894 = 11'h34d == cnt[10:0] ? $signed(-32'shf669) : $signed(_GEN_2893); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2895 = 11'h34e == cnt[10:0] ? $signed(-32'shf684) : $signed(_GEN_2894); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2896 = 11'h34f == cnt[10:0] ? $signed(-32'shf69f) : $signed(_GEN_2895); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2897 = 11'h350 == cnt[10:0] ? $signed(-32'shf6ba) : $signed(_GEN_2896); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2898 = 11'h351 == cnt[10:0] ? $signed(-32'shf6d5) : $signed(_GEN_2897); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2899 = 11'h352 == cnt[10:0] ? $signed(-32'shf6ef) : $signed(_GEN_2898); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2900 = 11'h353 == cnt[10:0] ? $signed(-32'shf70a) : $signed(_GEN_2899); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2901 = 11'h354 == cnt[10:0] ? $signed(-32'shf724) : $signed(_GEN_2900); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2902 = 11'h355 == cnt[10:0] ? $signed(-32'shf73e) : $signed(_GEN_2901); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2903 = 11'h356 == cnt[10:0] ? $signed(-32'shf758) : $signed(_GEN_2902); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2904 = 11'h357 == cnt[10:0] ? $signed(-32'shf772) : $signed(_GEN_2903); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2905 = 11'h358 == cnt[10:0] ? $signed(-32'shf78c) : $signed(_GEN_2904); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2906 = 11'h359 == cnt[10:0] ? $signed(-32'shf7a5) : $signed(_GEN_2905); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2907 = 11'h35a == cnt[10:0] ? $signed(-32'shf7bf) : $signed(_GEN_2906); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2908 = 11'h35b == cnt[10:0] ? $signed(-32'shf7d8) : $signed(_GEN_2907); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2909 = 11'h35c == cnt[10:0] ? $signed(-32'shf7f1) : $signed(_GEN_2908); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2910 = 11'h35d == cnt[10:0] ? $signed(-32'shf80a) : $signed(_GEN_2909); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2911 = 11'h35e == cnt[10:0] ? $signed(-32'shf823) : $signed(_GEN_2910); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2912 = 11'h35f == cnt[10:0] ? $signed(-32'shf83b) : $signed(_GEN_2911); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2913 = 11'h360 == cnt[10:0] ? $signed(-32'shf854) : $signed(_GEN_2912); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2914 = 11'h361 == cnt[10:0] ? $signed(-32'shf86c) : $signed(_GEN_2913); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2915 = 11'h362 == cnt[10:0] ? $signed(-32'shf885) : $signed(_GEN_2914); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2916 = 11'h363 == cnt[10:0] ? $signed(-32'shf89d) : $signed(_GEN_2915); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2917 = 11'h364 == cnt[10:0] ? $signed(-32'shf8b4) : $signed(_GEN_2916); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2918 = 11'h365 == cnt[10:0] ? $signed(-32'shf8cc) : $signed(_GEN_2917); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2919 = 11'h366 == cnt[10:0] ? $signed(-32'shf8e4) : $signed(_GEN_2918); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2920 = 11'h367 == cnt[10:0] ? $signed(-32'shf8fb) : $signed(_GEN_2919); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2921 = 11'h368 == cnt[10:0] ? $signed(-32'shf913) : $signed(_GEN_2920); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2922 = 11'h369 == cnt[10:0] ? $signed(-32'shf92a) : $signed(_GEN_2921); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2923 = 11'h36a == cnt[10:0] ? $signed(-32'shf941) : $signed(_GEN_2922); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2924 = 11'h36b == cnt[10:0] ? $signed(-32'shf958) : $signed(_GEN_2923); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2925 = 11'h36c == cnt[10:0] ? $signed(-32'shf96e) : $signed(_GEN_2924); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2926 = 11'h36d == cnt[10:0] ? $signed(-32'shf985) : $signed(_GEN_2925); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2927 = 11'h36e == cnt[10:0] ? $signed(-32'shf99b) : $signed(_GEN_2926); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2928 = 11'h36f == cnt[10:0] ? $signed(-32'shf9b2) : $signed(_GEN_2927); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2929 = 11'h370 == cnt[10:0] ? $signed(-32'shf9c8) : $signed(_GEN_2928); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2930 = 11'h371 == cnt[10:0] ? $signed(-32'shf9de) : $signed(_GEN_2929); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2931 = 11'h372 == cnt[10:0] ? $signed(-32'shf9f3) : $signed(_GEN_2930); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2932 = 11'h373 == cnt[10:0] ? $signed(-32'shfa09) : $signed(_GEN_2931); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2933 = 11'h374 == cnt[10:0] ? $signed(-32'shfa1f) : $signed(_GEN_2932); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2934 = 11'h375 == cnt[10:0] ? $signed(-32'shfa34) : $signed(_GEN_2933); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2935 = 11'h376 == cnt[10:0] ? $signed(-32'shfa49) : $signed(_GEN_2934); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2936 = 11'h377 == cnt[10:0] ? $signed(-32'shfa5e) : $signed(_GEN_2935); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2937 = 11'h378 == cnt[10:0] ? $signed(-32'shfa73) : $signed(_GEN_2936); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2938 = 11'h379 == cnt[10:0] ? $signed(-32'shfa88) : $signed(_GEN_2937); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2939 = 11'h37a == cnt[10:0] ? $signed(-32'shfa9c) : $signed(_GEN_2938); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2940 = 11'h37b == cnt[10:0] ? $signed(-32'shfab1) : $signed(_GEN_2939); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2941 = 11'h37c == cnt[10:0] ? $signed(-32'shfac5) : $signed(_GEN_2940); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2942 = 11'h37d == cnt[10:0] ? $signed(-32'shfad9) : $signed(_GEN_2941); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2943 = 11'h37e == cnt[10:0] ? $signed(-32'shfaed) : $signed(_GEN_2942); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2944 = 11'h37f == cnt[10:0] ? $signed(-32'shfb01) : $signed(_GEN_2943); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2945 = 11'h380 == cnt[10:0] ? $signed(-32'shfb15) : $signed(_GEN_2944); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2946 = 11'h381 == cnt[10:0] ? $signed(-32'shfb28) : $signed(_GEN_2945); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2947 = 11'h382 == cnt[10:0] ? $signed(-32'shfb3c) : $signed(_GEN_2946); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2948 = 11'h383 == cnt[10:0] ? $signed(-32'shfb4f) : $signed(_GEN_2947); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2949 = 11'h384 == cnt[10:0] ? $signed(-32'shfb62) : $signed(_GEN_2948); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2950 = 11'h385 == cnt[10:0] ? $signed(-32'shfb75) : $signed(_GEN_2949); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2951 = 11'h386 == cnt[10:0] ? $signed(-32'shfb88) : $signed(_GEN_2950); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2952 = 11'h387 == cnt[10:0] ? $signed(-32'shfb9a) : $signed(_GEN_2951); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2953 = 11'h388 == cnt[10:0] ? $signed(-32'shfbad) : $signed(_GEN_2952); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2954 = 11'h389 == cnt[10:0] ? $signed(-32'shfbbf) : $signed(_GEN_2953); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2955 = 11'h38a == cnt[10:0] ? $signed(-32'shfbd1) : $signed(_GEN_2954); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2956 = 11'h38b == cnt[10:0] ? $signed(-32'shfbe3) : $signed(_GEN_2955); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2957 = 11'h38c == cnt[10:0] ? $signed(-32'shfbf5) : $signed(_GEN_2956); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2958 = 11'h38d == cnt[10:0] ? $signed(-32'shfc07) : $signed(_GEN_2957); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2959 = 11'h38e == cnt[10:0] ? $signed(-32'shfc18) : $signed(_GEN_2958); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2960 = 11'h38f == cnt[10:0] ? $signed(-32'shfc2a) : $signed(_GEN_2959); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2961 = 11'h390 == cnt[10:0] ? $signed(-32'shfc3b) : $signed(_GEN_2960); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2962 = 11'h391 == cnt[10:0] ? $signed(-32'shfc4c) : $signed(_GEN_2961); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2963 = 11'h392 == cnt[10:0] ? $signed(-32'shfc5d) : $signed(_GEN_2962); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2964 = 11'h393 == cnt[10:0] ? $signed(-32'shfc6e) : $signed(_GEN_2963); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2965 = 11'h394 == cnt[10:0] ? $signed(-32'shfc7f) : $signed(_GEN_2964); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2966 = 11'h395 == cnt[10:0] ? $signed(-32'shfc8f) : $signed(_GEN_2965); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2967 = 11'h396 == cnt[10:0] ? $signed(-32'shfca0) : $signed(_GEN_2966); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2968 = 11'h397 == cnt[10:0] ? $signed(-32'shfcb0) : $signed(_GEN_2967); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2969 = 11'h398 == cnt[10:0] ? $signed(-32'shfcc0) : $signed(_GEN_2968); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2970 = 11'h399 == cnt[10:0] ? $signed(-32'shfcd0) : $signed(_GEN_2969); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2971 = 11'h39a == cnt[10:0] ? $signed(-32'shfcdf) : $signed(_GEN_2970); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2972 = 11'h39b == cnt[10:0] ? $signed(-32'shfcef) : $signed(_GEN_2971); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2973 = 11'h39c == cnt[10:0] ? $signed(-32'shfcfe) : $signed(_GEN_2972); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2974 = 11'h39d == cnt[10:0] ? $signed(-32'shfd0e) : $signed(_GEN_2973); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2975 = 11'h39e == cnt[10:0] ? $signed(-32'shfd1d) : $signed(_GEN_2974); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2976 = 11'h39f == cnt[10:0] ? $signed(-32'shfd2c) : $signed(_GEN_2975); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2977 = 11'h3a0 == cnt[10:0] ? $signed(-32'shfd3b) : $signed(_GEN_2976); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2978 = 11'h3a1 == cnt[10:0] ? $signed(-32'shfd49) : $signed(_GEN_2977); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2979 = 11'h3a2 == cnt[10:0] ? $signed(-32'shfd58) : $signed(_GEN_2978); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2980 = 11'h3a3 == cnt[10:0] ? $signed(-32'shfd66) : $signed(_GEN_2979); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2981 = 11'h3a4 == cnt[10:0] ? $signed(-32'shfd74) : $signed(_GEN_2980); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2982 = 11'h3a5 == cnt[10:0] ? $signed(-32'shfd83) : $signed(_GEN_2981); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2983 = 11'h3a6 == cnt[10:0] ? $signed(-32'shfd90) : $signed(_GEN_2982); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2984 = 11'h3a7 == cnt[10:0] ? $signed(-32'shfd9e) : $signed(_GEN_2983); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2985 = 11'h3a8 == cnt[10:0] ? $signed(-32'shfdac) : $signed(_GEN_2984); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2986 = 11'h3a9 == cnt[10:0] ? $signed(-32'shfdb9) : $signed(_GEN_2985); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2987 = 11'h3aa == cnt[10:0] ? $signed(-32'shfdc7) : $signed(_GEN_2986); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2988 = 11'h3ab == cnt[10:0] ? $signed(-32'shfdd4) : $signed(_GEN_2987); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2989 = 11'h3ac == cnt[10:0] ? $signed(-32'shfde1) : $signed(_GEN_2988); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2990 = 11'h3ad == cnt[10:0] ? $signed(-32'shfdee) : $signed(_GEN_2989); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2991 = 11'h3ae == cnt[10:0] ? $signed(-32'shfdfa) : $signed(_GEN_2990); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2992 = 11'h3af == cnt[10:0] ? $signed(-32'shfe07) : $signed(_GEN_2991); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2993 = 11'h3b0 == cnt[10:0] ? $signed(-32'shfe13) : $signed(_GEN_2992); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2994 = 11'h3b1 == cnt[10:0] ? $signed(-32'shfe1f) : $signed(_GEN_2993); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2995 = 11'h3b2 == cnt[10:0] ? $signed(-32'shfe2b) : $signed(_GEN_2994); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2996 = 11'h3b3 == cnt[10:0] ? $signed(-32'shfe37) : $signed(_GEN_2995); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2997 = 11'h3b4 == cnt[10:0] ? $signed(-32'shfe43) : $signed(_GEN_2996); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2998 = 11'h3b5 == cnt[10:0] ? $signed(-32'shfe4f) : $signed(_GEN_2997); // @[FFT.scala 35:12]
  wire [31:0] _GEN_2999 = 11'h3b6 == cnt[10:0] ? $signed(-32'shfe5a) : $signed(_GEN_2998); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3000 = 11'h3b7 == cnt[10:0] ? $signed(-32'shfe66) : $signed(_GEN_2999); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3001 = 11'h3b8 == cnt[10:0] ? $signed(-32'shfe71) : $signed(_GEN_3000); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3002 = 11'h3b9 == cnt[10:0] ? $signed(-32'shfe7c) : $signed(_GEN_3001); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3003 = 11'h3ba == cnt[10:0] ? $signed(-32'shfe87) : $signed(_GEN_3002); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3004 = 11'h3bb == cnt[10:0] ? $signed(-32'shfe91) : $signed(_GEN_3003); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3005 = 11'h3bc == cnt[10:0] ? $signed(-32'shfe9c) : $signed(_GEN_3004); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3006 = 11'h3bd == cnt[10:0] ? $signed(-32'shfea6) : $signed(_GEN_3005); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3007 = 11'h3be == cnt[10:0] ? $signed(-32'shfeb0) : $signed(_GEN_3006); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3008 = 11'h3bf == cnt[10:0] ? $signed(-32'shfeba) : $signed(_GEN_3007); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3009 = 11'h3c0 == cnt[10:0] ? $signed(-32'shfec4) : $signed(_GEN_3008); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3010 = 11'h3c1 == cnt[10:0] ? $signed(-32'shfece) : $signed(_GEN_3009); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3011 = 11'h3c2 == cnt[10:0] ? $signed(-32'shfed8) : $signed(_GEN_3010); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3012 = 11'h3c3 == cnt[10:0] ? $signed(-32'shfee1) : $signed(_GEN_3011); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3013 = 11'h3c4 == cnt[10:0] ? $signed(-32'shfeeb) : $signed(_GEN_3012); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3014 = 11'h3c5 == cnt[10:0] ? $signed(-32'shfef4) : $signed(_GEN_3013); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3015 = 11'h3c6 == cnt[10:0] ? $signed(-32'shfefd) : $signed(_GEN_3014); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3016 = 11'h3c7 == cnt[10:0] ? $signed(-32'shff06) : $signed(_GEN_3015); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3017 = 11'h3c8 == cnt[10:0] ? $signed(-32'shff0e) : $signed(_GEN_3016); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3018 = 11'h3c9 == cnt[10:0] ? $signed(-32'shff17) : $signed(_GEN_3017); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3019 = 11'h3ca == cnt[10:0] ? $signed(-32'shff1f) : $signed(_GEN_3018); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3020 = 11'h3cb == cnt[10:0] ? $signed(-32'shff28) : $signed(_GEN_3019); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3021 = 11'h3cc == cnt[10:0] ? $signed(-32'shff30) : $signed(_GEN_3020); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3022 = 11'h3cd == cnt[10:0] ? $signed(-32'shff38) : $signed(_GEN_3021); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3023 = 11'h3ce == cnt[10:0] ? $signed(-32'shff3f) : $signed(_GEN_3022); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3024 = 11'h3cf == cnt[10:0] ? $signed(-32'shff47) : $signed(_GEN_3023); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3025 = 11'h3d0 == cnt[10:0] ? $signed(-32'shff4e) : $signed(_GEN_3024); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3026 = 11'h3d1 == cnt[10:0] ? $signed(-32'shff56) : $signed(_GEN_3025); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3027 = 11'h3d2 == cnt[10:0] ? $signed(-32'shff5d) : $signed(_GEN_3026); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3028 = 11'h3d3 == cnt[10:0] ? $signed(-32'shff64) : $signed(_GEN_3027); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3029 = 11'h3d4 == cnt[10:0] ? $signed(-32'shff6b) : $signed(_GEN_3028); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3030 = 11'h3d5 == cnt[10:0] ? $signed(-32'shff71) : $signed(_GEN_3029); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3031 = 11'h3d6 == cnt[10:0] ? $signed(-32'shff78) : $signed(_GEN_3030); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3032 = 11'h3d7 == cnt[10:0] ? $signed(-32'shff7e) : $signed(_GEN_3031); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3033 = 11'h3d8 == cnt[10:0] ? $signed(-32'shff85) : $signed(_GEN_3032); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3034 = 11'h3d9 == cnt[10:0] ? $signed(-32'shff8b) : $signed(_GEN_3033); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3035 = 11'h3da == cnt[10:0] ? $signed(-32'shff91) : $signed(_GEN_3034); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3036 = 11'h3db == cnt[10:0] ? $signed(-32'shff96) : $signed(_GEN_3035); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3037 = 11'h3dc == cnt[10:0] ? $signed(-32'shff9c) : $signed(_GEN_3036); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3038 = 11'h3dd == cnt[10:0] ? $signed(-32'shffa2) : $signed(_GEN_3037); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3039 = 11'h3de == cnt[10:0] ? $signed(-32'shffa7) : $signed(_GEN_3038); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3040 = 11'h3df == cnt[10:0] ? $signed(-32'shffac) : $signed(_GEN_3039); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3041 = 11'h3e0 == cnt[10:0] ? $signed(-32'shffb1) : $signed(_GEN_3040); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3042 = 11'h3e1 == cnt[10:0] ? $signed(-32'shffb6) : $signed(_GEN_3041); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3043 = 11'h3e2 == cnt[10:0] ? $signed(-32'shffbb) : $signed(_GEN_3042); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3044 = 11'h3e3 == cnt[10:0] ? $signed(-32'shffbf) : $signed(_GEN_3043); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3045 = 11'h3e4 == cnt[10:0] ? $signed(-32'shffc4) : $signed(_GEN_3044); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3046 = 11'h3e5 == cnt[10:0] ? $signed(-32'shffc8) : $signed(_GEN_3045); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3047 = 11'h3e6 == cnt[10:0] ? $signed(-32'shffcc) : $signed(_GEN_3046); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3048 = 11'h3e7 == cnt[10:0] ? $signed(-32'shffd0) : $signed(_GEN_3047); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3049 = 11'h3e8 == cnt[10:0] ? $signed(-32'shffd4) : $signed(_GEN_3048); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3050 = 11'h3e9 == cnt[10:0] ? $signed(-32'shffd7) : $signed(_GEN_3049); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3051 = 11'h3ea == cnt[10:0] ? $signed(-32'shffdb) : $signed(_GEN_3050); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3052 = 11'h3eb == cnt[10:0] ? $signed(-32'shffde) : $signed(_GEN_3051); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3053 = 11'h3ec == cnt[10:0] ? $signed(-32'shffe1) : $signed(_GEN_3052); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3054 = 11'h3ed == cnt[10:0] ? $signed(-32'shffe4) : $signed(_GEN_3053); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3055 = 11'h3ee == cnt[10:0] ? $signed(-32'shffe7) : $signed(_GEN_3054); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3056 = 11'h3ef == cnt[10:0] ? $signed(-32'shffea) : $signed(_GEN_3055); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3057 = 11'h3f0 == cnt[10:0] ? $signed(-32'shffec) : $signed(_GEN_3056); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3058 = 11'h3f1 == cnt[10:0] ? $signed(-32'shffef) : $signed(_GEN_3057); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3059 = 11'h3f2 == cnt[10:0] ? $signed(-32'shfff1) : $signed(_GEN_3058); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3060 = 11'h3f3 == cnt[10:0] ? $signed(-32'shfff3) : $signed(_GEN_3059); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3061 = 11'h3f4 == cnt[10:0] ? $signed(-32'shfff5) : $signed(_GEN_3060); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3062 = 11'h3f5 == cnt[10:0] ? $signed(-32'shfff7) : $signed(_GEN_3061); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3063 = 11'h3f6 == cnt[10:0] ? $signed(-32'shfff8) : $signed(_GEN_3062); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3064 = 11'h3f7 == cnt[10:0] ? $signed(-32'shfffa) : $signed(_GEN_3063); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3065 = 11'h3f8 == cnt[10:0] ? $signed(-32'shfffb) : $signed(_GEN_3064); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3066 = 11'h3f9 == cnt[10:0] ? $signed(-32'shfffc) : $signed(_GEN_3065); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3067 = 11'h3fa == cnt[10:0] ? $signed(-32'shfffd) : $signed(_GEN_3066); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3068 = 11'h3fb == cnt[10:0] ? $signed(-32'shfffe) : $signed(_GEN_3067); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3069 = 11'h3fc == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_3068); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3070 = 11'h3fd == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_3069); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3071 = 11'h3fe == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_3070); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3072 = 11'h3ff == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_3071); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3073 = 11'h400 == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_3072); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3074 = 11'h401 == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_3073); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3075 = 11'h402 == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_3074); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3076 = 11'h403 == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_3075); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3077 = 11'h404 == cnt[10:0] ? $signed(-32'shffff) : $signed(_GEN_3076); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3078 = 11'h405 == cnt[10:0] ? $signed(-32'shfffe) : $signed(_GEN_3077); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3079 = 11'h406 == cnt[10:0] ? $signed(-32'shfffd) : $signed(_GEN_3078); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3080 = 11'h407 == cnt[10:0] ? $signed(-32'shfffc) : $signed(_GEN_3079); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3081 = 11'h408 == cnt[10:0] ? $signed(-32'shfffb) : $signed(_GEN_3080); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3082 = 11'h409 == cnt[10:0] ? $signed(-32'shfffa) : $signed(_GEN_3081); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3083 = 11'h40a == cnt[10:0] ? $signed(-32'shfff8) : $signed(_GEN_3082); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3084 = 11'h40b == cnt[10:0] ? $signed(-32'shfff7) : $signed(_GEN_3083); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3085 = 11'h40c == cnt[10:0] ? $signed(-32'shfff5) : $signed(_GEN_3084); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3086 = 11'h40d == cnt[10:0] ? $signed(-32'shfff3) : $signed(_GEN_3085); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3087 = 11'h40e == cnt[10:0] ? $signed(-32'shfff1) : $signed(_GEN_3086); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3088 = 11'h40f == cnt[10:0] ? $signed(-32'shffef) : $signed(_GEN_3087); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3089 = 11'h410 == cnt[10:0] ? $signed(-32'shffec) : $signed(_GEN_3088); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3090 = 11'h411 == cnt[10:0] ? $signed(-32'shffea) : $signed(_GEN_3089); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3091 = 11'h412 == cnt[10:0] ? $signed(-32'shffe7) : $signed(_GEN_3090); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3092 = 11'h413 == cnt[10:0] ? $signed(-32'shffe4) : $signed(_GEN_3091); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3093 = 11'h414 == cnt[10:0] ? $signed(-32'shffe1) : $signed(_GEN_3092); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3094 = 11'h415 == cnt[10:0] ? $signed(-32'shffde) : $signed(_GEN_3093); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3095 = 11'h416 == cnt[10:0] ? $signed(-32'shffdb) : $signed(_GEN_3094); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3096 = 11'h417 == cnt[10:0] ? $signed(-32'shffd7) : $signed(_GEN_3095); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3097 = 11'h418 == cnt[10:0] ? $signed(-32'shffd4) : $signed(_GEN_3096); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3098 = 11'h419 == cnt[10:0] ? $signed(-32'shffd0) : $signed(_GEN_3097); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3099 = 11'h41a == cnt[10:0] ? $signed(-32'shffcc) : $signed(_GEN_3098); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3100 = 11'h41b == cnt[10:0] ? $signed(-32'shffc8) : $signed(_GEN_3099); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3101 = 11'h41c == cnt[10:0] ? $signed(-32'shffc4) : $signed(_GEN_3100); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3102 = 11'h41d == cnt[10:0] ? $signed(-32'shffbf) : $signed(_GEN_3101); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3103 = 11'h41e == cnt[10:0] ? $signed(-32'shffbb) : $signed(_GEN_3102); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3104 = 11'h41f == cnt[10:0] ? $signed(-32'shffb6) : $signed(_GEN_3103); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3105 = 11'h420 == cnt[10:0] ? $signed(-32'shffb1) : $signed(_GEN_3104); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3106 = 11'h421 == cnt[10:0] ? $signed(-32'shffac) : $signed(_GEN_3105); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3107 = 11'h422 == cnt[10:0] ? $signed(-32'shffa7) : $signed(_GEN_3106); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3108 = 11'h423 == cnt[10:0] ? $signed(-32'shffa2) : $signed(_GEN_3107); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3109 = 11'h424 == cnt[10:0] ? $signed(-32'shff9c) : $signed(_GEN_3108); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3110 = 11'h425 == cnt[10:0] ? $signed(-32'shff96) : $signed(_GEN_3109); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3111 = 11'h426 == cnt[10:0] ? $signed(-32'shff91) : $signed(_GEN_3110); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3112 = 11'h427 == cnt[10:0] ? $signed(-32'shff8b) : $signed(_GEN_3111); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3113 = 11'h428 == cnt[10:0] ? $signed(-32'shff85) : $signed(_GEN_3112); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3114 = 11'h429 == cnt[10:0] ? $signed(-32'shff7e) : $signed(_GEN_3113); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3115 = 11'h42a == cnt[10:0] ? $signed(-32'shff78) : $signed(_GEN_3114); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3116 = 11'h42b == cnt[10:0] ? $signed(-32'shff71) : $signed(_GEN_3115); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3117 = 11'h42c == cnt[10:0] ? $signed(-32'shff6b) : $signed(_GEN_3116); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3118 = 11'h42d == cnt[10:0] ? $signed(-32'shff64) : $signed(_GEN_3117); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3119 = 11'h42e == cnt[10:0] ? $signed(-32'shff5d) : $signed(_GEN_3118); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3120 = 11'h42f == cnt[10:0] ? $signed(-32'shff56) : $signed(_GEN_3119); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3121 = 11'h430 == cnt[10:0] ? $signed(-32'shff4e) : $signed(_GEN_3120); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3122 = 11'h431 == cnt[10:0] ? $signed(-32'shff47) : $signed(_GEN_3121); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3123 = 11'h432 == cnt[10:0] ? $signed(-32'shff3f) : $signed(_GEN_3122); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3124 = 11'h433 == cnt[10:0] ? $signed(-32'shff38) : $signed(_GEN_3123); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3125 = 11'h434 == cnt[10:0] ? $signed(-32'shff30) : $signed(_GEN_3124); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3126 = 11'h435 == cnt[10:0] ? $signed(-32'shff28) : $signed(_GEN_3125); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3127 = 11'h436 == cnt[10:0] ? $signed(-32'shff1f) : $signed(_GEN_3126); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3128 = 11'h437 == cnt[10:0] ? $signed(-32'shff17) : $signed(_GEN_3127); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3129 = 11'h438 == cnt[10:0] ? $signed(-32'shff0e) : $signed(_GEN_3128); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3130 = 11'h439 == cnt[10:0] ? $signed(-32'shff06) : $signed(_GEN_3129); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3131 = 11'h43a == cnt[10:0] ? $signed(-32'shfefd) : $signed(_GEN_3130); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3132 = 11'h43b == cnt[10:0] ? $signed(-32'shfef4) : $signed(_GEN_3131); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3133 = 11'h43c == cnt[10:0] ? $signed(-32'shfeeb) : $signed(_GEN_3132); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3134 = 11'h43d == cnt[10:0] ? $signed(-32'shfee1) : $signed(_GEN_3133); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3135 = 11'h43e == cnt[10:0] ? $signed(-32'shfed8) : $signed(_GEN_3134); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3136 = 11'h43f == cnt[10:0] ? $signed(-32'shfece) : $signed(_GEN_3135); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3137 = 11'h440 == cnt[10:0] ? $signed(-32'shfec4) : $signed(_GEN_3136); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3138 = 11'h441 == cnt[10:0] ? $signed(-32'shfeba) : $signed(_GEN_3137); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3139 = 11'h442 == cnt[10:0] ? $signed(-32'shfeb0) : $signed(_GEN_3138); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3140 = 11'h443 == cnt[10:0] ? $signed(-32'shfea6) : $signed(_GEN_3139); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3141 = 11'h444 == cnt[10:0] ? $signed(-32'shfe9c) : $signed(_GEN_3140); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3142 = 11'h445 == cnt[10:0] ? $signed(-32'shfe91) : $signed(_GEN_3141); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3143 = 11'h446 == cnt[10:0] ? $signed(-32'shfe87) : $signed(_GEN_3142); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3144 = 11'h447 == cnt[10:0] ? $signed(-32'shfe7c) : $signed(_GEN_3143); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3145 = 11'h448 == cnt[10:0] ? $signed(-32'shfe71) : $signed(_GEN_3144); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3146 = 11'h449 == cnt[10:0] ? $signed(-32'shfe66) : $signed(_GEN_3145); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3147 = 11'h44a == cnt[10:0] ? $signed(-32'shfe5a) : $signed(_GEN_3146); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3148 = 11'h44b == cnt[10:0] ? $signed(-32'shfe4f) : $signed(_GEN_3147); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3149 = 11'h44c == cnt[10:0] ? $signed(-32'shfe43) : $signed(_GEN_3148); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3150 = 11'h44d == cnt[10:0] ? $signed(-32'shfe37) : $signed(_GEN_3149); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3151 = 11'h44e == cnt[10:0] ? $signed(-32'shfe2b) : $signed(_GEN_3150); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3152 = 11'h44f == cnt[10:0] ? $signed(-32'shfe1f) : $signed(_GEN_3151); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3153 = 11'h450 == cnt[10:0] ? $signed(-32'shfe13) : $signed(_GEN_3152); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3154 = 11'h451 == cnt[10:0] ? $signed(-32'shfe07) : $signed(_GEN_3153); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3155 = 11'h452 == cnt[10:0] ? $signed(-32'shfdfa) : $signed(_GEN_3154); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3156 = 11'h453 == cnt[10:0] ? $signed(-32'shfdee) : $signed(_GEN_3155); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3157 = 11'h454 == cnt[10:0] ? $signed(-32'shfde1) : $signed(_GEN_3156); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3158 = 11'h455 == cnt[10:0] ? $signed(-32'shfdd4) : $signed(_GEN_3157); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3159 = 11'h456 == cnt[10:0] ? $signed(-32'shfdc7) : $signed(_GEN_3158); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3160 = 11'h457 == cnt[10:0] ? $signed(-32'shfdb9) : $signed(_GEN_3159); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3161 = 11'h458 == cnt[10:0] ? $signed(-32'shfdac) : $signed(_GEN_3160); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3162 = 11'h459 == cnt[10:0] ? $signed(-32'shfd9e) : $signed(_GEN_3161); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3163 = 11'h45a == cnt[10:0] ? $signed(-32'shfd90) : $signed(_GEN_3162); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3164 = 11'h45b == cnt[10:0] ? $signed(-32'shfd83) : $signed(_GEN_3163); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3165 = 11'h45c == cnt[10:0] ? $signed(-32'shfd74) : $signed(_GEN_3164); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3166 = 11'h45d == cnt[10:0] ? $signed(-32'shfd66) : $signed(_GEN_3165); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3167 = 11'h45e == cnt[10:0] ? $signed(-32'shfd58) : $signed(_GEN_3166); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3168 = 11'h45f == cnt[10:0] ? $signed(-32'shfd49) : $signed(_GEN_3167); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3169 = 11'h460 == cnt[10:0] ? $signed(-32'shfd3b) : $signed(_GEN_3168); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3170 = 11'h461 == cnt[10:0] ? $signed(-32'shfd2c) : $signed(_GEN_3169); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3171 = 11'h462 == cnt[10:0] ? $signed(-32'shfd1d) : $signed(_GEN_3170); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3172 = 11'h463 == cnt[10:0] ? $signed(-32'shfd0e) : $signed(_GEN_3171); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3173 = 11'h464 == cnt[10:0] ? $signed(-32'shfcfe) : $signed(_GEN_3172); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3174 = 11'h465 == cnt[10:0] ? $signed(-32'shfcef) : $signed(_GEN_3173); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3175 = 11'h466 == cnt[10:0] ? $signed(-32'shfcdf) : $signed(_GEN_3174); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3176 = 11'h467 == cnt[10:0] ? $signed(-32'shfcd0) : $signed(_GEN_3175); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3177 = 11'h468 == cnt[10:0] ? $signed(-32'shfcc0) : $signed(_GEN_3176); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3178 = 11'h469 == cnt[10:0] ? $signed(-32'shfcb0) : $signed(_GEN_3177); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3179 = 11'h46a == cnt[10:0] ? $signed(-32'shfca0) : $signed(_GEN_3178); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3180 = 11'h46b == cnt[10:0] ? $signed(-32'shfc8f) : $signed(_GEN_3179); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3181 = 11'h46c == cnt[10:0] ? $signed(-32'shfc7f) : $signed(_GEN_3180); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3182 = 11'h46d == cnt[10:0] ? $signed(-32'shfc6e) : $signed(_GEN_3181); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3183 = 11'h46e == cnt[10:0] ? $signed(-32'shfc5d) : $signed(_GEN_3182); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3184 = 11'h46f == cnt[10:0] ? $signed(-32'shfc4c) : $signed(_GEN_3183); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3185 = 11'h470 == cnt[10:0] ? $signed(-32'shfc3b) : $signed(_GEN_3184); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3186 = 11'h471 == cnt[10:0] ? $signed(-32'shfc2a) : $signed(_GEN_3185); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3187 = 11'h472 == cnt[10:0] ? $signed(-32'shfc18) : $signed(_GEN_3186); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3188 = 11'h473 == cnt[10:0] ? $signed(-32'shfc07) : $signed(_GEN_3187); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3189 = 11'h474 == cnt[10:0] ? $signed(-32'shfbf5) : $signed(_GEN_3188); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3190 = 11'h475 == cnt[10:0] ? $signed(-32'shfbe3) : $signed(_GEN_3189); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3191 = 11'h476 == cnt[10:0] ? $signed(-32'shfbd1) : $signed(_GEN_3190); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3192 = 11'h477 == cnt[10:0] ? $signed(-32'shfbbf) : $signed(_GEN_3191); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3193 = 11'h478 == cnt[10:0] ? $signed(-32'shfbad) : $signed(_GEN_3192); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3194 = 11'h479 == cnt[10:0] ? $signed(-32'shfb9a) : $signed(_GEN_3193); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3195 = 11'h47a == cnt[10:0] ? $signed(-32'shfb88) : $signed(_GEN_3194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3196 = 11'h47b == cnt[10:0] ? $signed(-32'shfb75) : $signed(_GEN_3195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3197 = 11'h47c == cnt[10:0] ? $signed(-32'shfb62) : $signed(_GEN_3196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3198 = 11'h47d == cnt[10:0] ? $signed(-32'shfb4f) : $signed(_GEN_3197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3199 = 11'h47e == cnt[10:0] ? $signed(-32'shfb3c) : $signed(_GEN_3198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3200 = 11'h47f == cnt[10:0] ? $signed(-32'shfb28) : $signed(_GEN_3199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3201 = 11'h480 == cnt[10:0] ? $signed(-32'shfb15) : $signed(_GEN_3200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3202 = 11'h481 == cnt[10:0] ? $signed(-32'shfb01) : $signed(_GEN_3201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3203 = 11'h482 == cnt[10:0] ? $signed(-32'shfaed) : $signed(_GEN_3202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3204 = 11'h483 == cnt[10:0] ? $signed(-32'shfad9) : $signed(_GEN_3203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3205 = 11'h484 == cnt[10:0] ? $signed(-32'shfac5) : $signed(_GEN_3204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3206 = 11'h485 == cnt[10:0] ? $signed(-32'shfab1) : $signed(_GEN_3205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3207 = 11'h486 == cnt[10:0] ? $signed(-32'shfa9c) : $signed(_GEN_3206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3208 = 11'h487 == cnt[10:0] ? $signed(-32'shfa88) : $signed(_GEN_3207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3209 = 11'h488 == cnt[10:0] ? $signed(-32'shfa73) : $signed(_GEN_3208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3210 = 11'h489 == cnt[10:0] ? $signed(-32'shfa5e) : $signed(_GEN_3209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3211 = 11'h48a == cnt[10:0] ? $signed(-32'shfa49) : $signed(_GEN_3210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3212 = 11'h48b == cnt[10:0] ? $signed(-32'shfa34) : $signed(_GEN_3211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3213 = 11'h48c == cnt[10:0] ? $signed(-32'shfa1f) : $signed(_GEN_3212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3214 = 11'h48d == cnt[10:0] ? $signed(-32'shfa09) : $signed(_GEN_3213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3215 = 11'h48e == cnt[10:0] ? $signed(-32'shf9f3) : $signed(_GEN_3214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3216 = 11'h48f == cnt[10:0] ? $signed(-32'shf9de) : $signed(_GEN_3215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3217 = 11'h490 == cnt[10:0] ? $signed(-32'shf9c8) : $signed(_GEN_3216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3218 = 11'h491 == cnt[10:0] ? $signed(-32'shf9b2) : $signed(_GEN_3217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3219 = 11'h492 == cnt[10:0] ? $signed(-32'shf99b) : $signed(_GEN_3218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3220 = 11'h493 == cnt[10:0] ? $signed(-32'shf985) : $signed(_GEN_3219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3221 = 11'h494 == cnt[10:0] ? $signed(-32'shf96e) : $signed(_GEN_3220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3222 = 11'h495 == cnt[10:0] ? $signed(-32'shf958) : $signed(_GEN_3221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3223 = 11'h496 == cnt[10:0] ? $signed(-32'shf941) : $signed(_GEN_3222); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3224 = 11'h497 == cnt[10:0] ? $signed(-32'shf92a) : $signed(_GEN_3223); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3225 = 11'h498 == cnt[10:0] ? $signed(-32'shf913) : $signed(_GEN_3224); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3226 = 11'h499 == cnt[10:0] ? $signed(-32'shf8fb) : $signed(_GEN_3225); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3227 = 11'h49a == cnt[10:0] ? $signed(-32'shf8e4) : $signed(_GEN_3226); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3228 = 11'h49b == cnt[10:0] ? $signed(-32'shf8cc) : $signed(_GEN_3227); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3229 = 11'h49c == cnt[10:0] ? $signed(-32'shf8b4) : $signed(_GEN_3228); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3230 = 11'h49d == cnt[10:0] ? $signed(-32'shf89d) : $signed(_GEN_3229); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3231 = 11'h49e == cnt[10:0] ? $signed(-32'shf885) : $signed(_GEN_3230); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3232 = 11'h49f == cnt[10:0] ? $signed(-32'shf86c) : $signed(_GEN_3231); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3233 = 11'h4a0 == cnt[10:0] ? $signed(-32'shf854) : $signed(_GEN_3232); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3234 = 11'h4a1 == cnt[10:0] ? $signed(-32'shf83b) : $signed(_GEN_3233); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3235 = 11'h4a2 == cnt[10:0] ? $signed(-32'shf823) : $signed(_GEN_3234); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3236 = 11'h4a3 == cnt[10:0] ? $signed(-32'shf80a) : $signed(_GEN_3235); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3237 = 11'h4a4 == cnt[10:0] ? $signed(-32'shf7f1) : $signed(_GEN_3236); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3238 = 11'h4a5 == cnt[10:0] ? $signed(-32'shf7d8) : $signed(_GEN_3237); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3239 = 11'h4a6 == cnt[10:0] ? $signed(-32'shf7bf) : $signed(_GEN_3238); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3240 = 11'h4a7 == cnt[10:0] ? $signed(-32'shf7a5) : $signed(_GEN_3239); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3241 = 11'h4a8 == cnt[10:0] ? $signed(-32'shf78c) : $signed(_GEN_3240); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3242 = 11'h4a9 == cnt[10:0] ? $signed(-32'shf772) : $signed(_GEN_3241); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3243 = 11'h4aa == cnt[10:0] ? $signed(-32'shf758) : $signed(_GEN_3242); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3244 = 11'h4ab == cnt[10:0] ? $signed(-32'shf73e) : $signed(_GEN_3243); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3245 = 11'h4ac == cnt[10:0] ? $signed(-32'shf724) : $signed(_GEN_3244); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3246 = 11'h4ad == cnt[10:0] ? $signed(-32'shf70a) : $signed(_GEN_3245); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3247 = 11'h4ae == cnt[10:0] ? $signed(-32'shf6ef) : $signed(_GEN_3246); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3248 = 11'h4af == cnt[10:0] ? $signed(-32'shf6d5) : $signed(_GEN_3247); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3249 = 11'h4b0 == cnt[10:0] ? $signed(-32'shf6ba) : $signed(_GEN_3248); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3250 = 11'h4b1 == cnt[10:0] ? $signed(-32'shf69f) : $signed(_GEN_3249); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3251 = 11'h4b2 == cnt[10:0] ? $signed(-32'shf684) : $signed(_GEN_3250); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3252 = 11'h4b3 == cnt[10:0] ? $signed(-32'shf669) : $signed(_GEN_3251); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3253 = 11'h4b4 == cnt[10:0] ? $signed(-32'shf64e) : $signed(_GEN_3252); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3254 = 11'h4b5 == cnt[10:0] ? $signed(-32'shf632) : $signed(_GEN_3253); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3255 = 11'h4b6 == cnt[10:0] ? $signed(-32'shf616) : $signed(_GEN_3254); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3256 = 11'h4b7 == cnt[10:0] ? $signed(-32'shf5fb) : $signed(_GEN_3255); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3257 = 11'h4b8 == cnt[10:0] ? $signed(-32'shf5df) : $signed(_GEN_3256); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3258 = 11'h4b9 == cnt[10:0] ? $signed(-32'shf5c3) : $signed(_GEN_3257); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3259 = 11'h4ba == cnt[10:0] ? $signed(-32'shf5a6) : $signed(_GEN_3258); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3260 = 11'h4bb == cnt[10:0] ? $signed(-32'shf58a) : $signed(_GEN_3259); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3261 = 11'h4bc == cnt[10:0] ? $signed(-32'shf56e) : $signed(_GEN_3260); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3262 = 11'h4bd == cnt[10:0] ? $signed(-32'shf551) : $signed(_GEN_3261); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3263 = 11'h4be == cnt[10:0] ? $signed(-32'shf534) : $signed(_GEN_3262); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3264 = 11'h4bf == cnt[10:0] ? $signed(-32'shf517) : $signed(_GEN_3263); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3265 = 11'h4c0 == cnt[10:0] ? $signed(-32'shf4fa) : $signed(_GEN_3264); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3266 = 11'h4c1 == cnt[10:0] ? $signed(-32'shf4dd) : $signed(_GEN_3265); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3267 = 11'h4c2 == cnt[10:0] ? $signed(-32'shf4bf) : $signed(_GEN_3266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3268 = 11'h4c3 == cnt[10:0] ? $signed(-32'shf4a2) : $signed(_GEN_3267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3269 = 11'h4c4 == cnt[10:0] ? $signed(-32'shf484) : $signed(_GEN_3268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3270 = 11'h4c5 == cnt[10:0] ? $signed(-32'shf466) : $signed(_GEN_3269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3271 = 11'h4c6 == cnt[10:0] ? $signed(-32'shf448) : $signed(_GEN_3270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3272 = 11'h4c7 == cnt[10:0] ? $signed(-32'shf42a) : $signed(_GEN_3271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3273 = 11'h4c8 == cnt[10:0] ? $signed(-32'shf40c) : $signed(_GEN_3272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3274 = 11'h4c9 == cnt[10:0] ? $signed(-32'shf3ed) : $signed(_GEN_3273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3275 = 11'h4ca == cnt[10:0] ? $signed(-32'shf3cf) : $signed(_GEN_3274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3276 = 11'h4cb == cnt[10:0] ? $signed(-32'shf3b0) : $signed(_GEN_3275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3277 = 11'h4cc == cnt[10:0] ? $signed(-32'shf391) : $signed(_GEN_3276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3278 = 11'h4cd == cnt[10:0] ? $signed(-32'shf372) : $signed(_GEN_3277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3279 = 11'h4ce == cnt[10:0] ? $signed(-32'shf353) : $signed(_GEN_3278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3280 = 11'h4cf == cnt[10:0] ? $signed(-32'shf334) : $signed(_GEN_3279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3281 = 11'h4d0 == cnt[10:0] ? $signed(-32'shf314) : $signed(_GEN_3280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3282 = 11'h4d1 == cnt[10:0] ? $signed(-32'shf2f5) : $signed(_GEN_3281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3283 = 11'h4d2 == cnt[10:0] ? $signed(-32'shf2d5) : $signed(_GEN_3282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3284 = 11'h4d3 == cnt[10:0] ? $signed(-32'shf2b5) : $signed(_GEN_3283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3285 = 11'h4d4 == cnt[10:0] ? $signed(-32'shf295) : $signed(_GEN_3284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3286 = 11'h4d5 == cnt[10:0] ? $signed(-32'shf275) : $signed(_GEN_3285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3287 = 11'h4d6 == cnt[10:0] ? $signed(-32'shf254) : $signed(_GEN_3286); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3288 = 11'h4d7 == cnt[10:0] ? $signed(-32'shf234) : $signed(_GEN_3287); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3289 = 11'h4d8 == cnt[10:0] ? $signed(-32'shf213) : $signed(_GEN_3288); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3290 = 11'h4d9 == cnt[10:0] ? $signed(-32'shf1f3) : $signed(_GEN_3289); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3291 = 11'h4da == cnt[10:0] ? $signed(-32'shf1d2) : $signed(_GEN_3290); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3292 = 11'h4db == cnt[10:0] ? $signed(-32'shf1b1) : $signed(_GEN_3291); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3293 = 11'h4dc == cnt[10:0] ? $signed(-32'shf18f) : $signed(_GEN_3292); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3294 = 11'h4dd == cnt[10:0] ? $signed(-32'shf16e) : $signed(_GEN_3293); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3295 = 11'h4de == cnt[10:0] ? $signed(-32'shf14c) : $signed(_GEN_3294); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3296 = 11'h4df == cnt[10:0] ? $signed(-32'shf12b) : $signed(_GEN_3295); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3297 = 11'h4e0 == cnt[10:0] ? $signed(-32'shf109) : $signed(_GEN_3296); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3298 = 11'h4e1 == cnt[10:0] ? $signed(-32'shf0e7) : $signed(_GEN_3297); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3299 = 11'h4e2 == cnt[10:0] ? $signed(-32'shf0c5) : $signed(_GEN_3298); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3300 = 11'h4e3 == cnt[10:0] ? $signed(-32'shf0a3) : $signed(_GEN_3299); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3301 = 11'h4e4 == cnt[10:0] ? $signed(-32'shf080) : $signed(_GEN_3300); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3302 = 11'h4e5 == cnt[10:0] ? $signed(-32'shf05e) : $signed(_GEN_3301); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3303 = 11'h4e6 == cnt[10:0] ? $signed(-32'shf03b) : $signed(_GEN_3302); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3304 = 11'h4e7 == cnt[10:0] ? $signed(-32'shf018) : $signed(_GEN_3303); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3305 = 11'h4e8 == cnt[10:0] ? $signed(-32'sheff5) : $signed(_GEN_3304); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3306 = 11'h4e9 == cnt[10:0] ? $signed(-32'shefd2) : $signed(_GEN_3305); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3307 = 11'h4ea == cnt[10:0] ? $signed(-32'shefaf) : $signed(_GEN_3306); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3308 = 11'h4eb == cnt[10:0] ? $signed(-32'shef8c) : $signed(_GEN_3307); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3309 = 11'h4ec == cnt[10:0] ? $signed(-32'shef68) : $signed(_GEN_3308); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3310 = 11'h4ed == cnt[10:0] ? $signed(-32'shef45) : $signed(_GEN_3309); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3311 = 11'h4ee == cnt[10:0] ? $signed(-32'shef21) : $signed(_GEN_3310); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3312 = 11'h4ef == cnt[10:0] ? $signed(-32'sheefd) : $signed(_GEN_3311); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3313 = 11'h4f0 == cnt[10:0] ? $signed(-32'sheed9) : $signed(_GEN_3312); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3314 = 11'h4f1 == cnt[10:0] ? $signed(-32'sheeb4) : $signed(_GEN_3313); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3315 = 11'h4f2 == cnt[10:0] ? $signed(-32'shee90) : $signed(_GEN_3314); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3316 = 11'h4f3 == cnt[10:0] ? $signed(-32'shee6b) : $signed(_GEN_3315); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3317 = 11'h4f4 == cnt[10:0] ? $signed(-32'shee47) : $signed(_GEN_3316); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3318 = 11'h4f5 == cnt[10:0] ? $signed(-32'shee22) : $signed(_GEN_3317); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3319 = 11'h4f6 == cnt[10:0] ? $signed(-32'shedfd) : $signed(_GEN_3318); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3320 = 11'h4f7 == cnt[10:0] ? $signed(-32'shedd8) : $signed(_GEN_3319); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3321 = 11'h4f8 == cnt[10:0] ? $signed(-32'shedb3) : $signed(_GEN_3320); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3322 = 11'h4f9 == cnt[10:0] ? $signed(-32'shed8d) : $signed(_GEN_3321); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3323 = 11'h4fa == cnt[10:0] ? $signed(-32'shed68) : $signed(_GEN_3322); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3324 = 11'h4fb == cnt[10:0] ? $signed(-32'shed42) : $signed(_GEN_3323); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3325 = 11'h4fc == cnt[10:0] ? $signed(-32'shed1c) : $signed(_GEN_3324); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3326 = 11'h4fd == cnt[10:0] ? $signed(-32'shecf6) : $signed(_GEN_3325); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3327 = 11'h4fe == cnt[10:0] ? $signed(-32'shecd0) : $signed(_GEN_3326); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3328 = 11'h4ff == cnt[10:0] ? $signed(-32'shecaa) : $signed(_GEN_3327); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3329 = 11'h500 == cnt[10:0] ? $signed(-32'shec83) : $signed(_GEN_3328); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3330 = 11'h501 == cnt[10:0] ? $signed(-32'shec5d) : $signed(_GEN_3329); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3331 = 11'h502 == cnt[10:0] ? $signed(-32'shec36) : $signed(_GEN_3330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3332 = 11'h503 == cnt[10:0] ? $signed(-32'shec0f) : $signed(_GEN_3331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3333 = 11'h504 == cnt[10:0] ? $signed(-32'shebe8) : $signed(_GEN_3332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3334 = 11'h505 == cnt[10:0] ? $signed(-32'shebc1) : $signed(_GEN_3333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3335 = 11'h506 == cnt[10:0] ? $signed(-32'sheb9a) : $signed(_GEN_3334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3336 = 11'h507 == cnt[10:0] ? $signed(-32'sheb73) : $signed(_GEN_3335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3337 = 11'h508 == cnt[10:0] ? $signed(-32'sheb4b) : $signed(_GEN_3336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3338 = 11'h509 == cnt[10:0] ? $signed(-32'sheb23) : $signed(_GEN_3337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3339 = 11'h50a == cnt[10:0] ? $signed(-32'sheafc) : $signed(_GEN_3338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3340 = 11'h50b == cnt[10:0] ? $signed(-32'shead4) : $signed(_GEN_3339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3341 = 11'h50c == cnt[10:0] ? $signed(-32'sheaab) : $signed(_GEN_3340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3342 = 11'h50d == cnt[10:0] ? $signed(-32'shea83) : $signed(_GEN_3341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3343 = 11'h50e == cnt[10:0] ? $signed(-32'shea5b) : $signed(_GEN_3342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3344 = 11'h50f == cnt[10:0] ? $signed(-32'shea32) : $signed(_GEN_3343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3345 = 11'h510 == cnt[10:0] ? $signed(-32'shea0a) : $signed(_GEN_3344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3346 = 11'h511 == cnt[10:0] ? $signed(-32'she9e1) : $signed(_GEN_3345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3347 = 11'h512 == cnt[10:0] ? $signed(-32'she9b8) : $signed(_GEN_3346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3348 = 11'h513 == cnt[10:0] ? $signed(-32'she98f) : $signed(_GEN_3347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3349 = 11'h514 == cnt[10:0] ? $signed(-32'she966) : $signed(_GEN_3348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3350 = 11'h515 == cnt[10:0] ? $signed(-32'she93c) : $signed(_GEN_3349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3351 = 11'h516 == cnt[10:0] ? $signed(-32'she913) : $signed(_GEN_3350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3352 = 11'h517 == cnt[10:0] ? $signed(-32'she8e9) : $signed(_GEN_3351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3353 = 11'h518 == cnt[10:0] ? $signed(-32'she8bf) : $signed(_GEN_3352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3354 = 11'h519 == cnt[10:0] ? $signed(-32'she895) : $signed(_GEN_3353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3355 = 11'h51a == cnt[10:0] ? $signed(-32'she86b) : $signed(_GEN_3354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3356 = 11'h51b == cnt[10:0] ? $signed(-32'she841) : $signed(_GEN_3355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3357 = 11'h51c == cnt[10:0] ? $signed(-32'she817) : $signed(_GEN_3356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3358 = 11'h51d == cnt[10:0] ? $signed(-32'she7ec) : $signed(_GEN_3357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3359 = 11'h51e == cnt[10:0] ? $signed(-32'she7c2) : $signed(_GEN_3358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3360 = 11'h51f == cnt[10:0] ? $signed(-32'she797) : $signed(_GEN_3359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3361 = 11'h520 == cnt[10:0] ? $signed(-32'she76c) : $signed(_GEN_3360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3362 = 11'h521 == cnt[10:0] ? $signed(-32'she741) : $signed(_GEN_3361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3363 = 11'h522 == cnt[10:0] ? $signed(-32'she716) : $signed(_GEN_3362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3364 = 11'h523 == cnt[10:0] ? $signed(-32'she6ea) : $signed(_GEN_3363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3365 = 11'h524 == cnt[10:0] ? $signed(-32'she6bf) : $signed(_GEN_3364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3366 = 11'h525 == cnt[10:0] ? $signed(-32'she693) : $signed(_GEN_3365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3367 = 11'h526 == cnt[10:0] ? $signed(-32'she667) : $signed(_GEN_3366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3368 = 11'h527 == cnt[10:0] ? $signed(-32'she63c) : $signed(_GEN_3367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3369 = 11'h528 == cnt[10:0] ? $signed(-32'she610) : $signed(_GEN_3368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3370 = 11'h529 == cnt[10:0] ? $signed(-32'she5e3) : $signed(_GEN_3369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3371 = 11'h52a == cnt[10:0] ? $signed(-32'she5b7) : $signed(_GEN_3370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3372 = 11'h52b == cnt[10:0] ? $signed(-32'she58b) : $signed(_GEN_3371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3373 = 11'h52c == cnt[10:0] ? $signed(-32'she55e) : $signed(_GEN_3372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3374 = 11'h52d == cnt[10:0] ? $signed(-32'she531) : $signed(_GEN_3373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3375 = 11'h52e == cnt[10:0] ? $signed(-32'she504) : $signed(_GEN_3374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3376 = 11'h52f == cnt[10:0] ? $signed(-32'she4d7) : $signed(_GEN_3375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3377 = 11'h530 == cnt[10:0] ? $signed(-32'she4aa) : $signed(_GEN_3376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3378 = 11'h531 == cnt[10:0] ? $signed(-32'she47d) : $signed(_GEN_3377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3379 = 11'h532 == cnt[10:0] ? $signed(-32'she450) : $signed(_GEN_3378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3380 = 11'h533 == cnt[10:0] ? $signed(-32'she422) : $signed(_GEN_3379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3381 = 11'h534 == cnt[10:0] ? $signed(-32'she3f4) : $signed(_GEN_3380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3382 = 11'h535 == cnt[10:0] ? $signed(-32'she3c7) : $signed(_GEN_3381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3383 = 11'h536 == cnt[10:0] ? $signed(-32'she399) : $signed(_GEN_3382); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3384 = 11'h537 == cnt[10:0] ? $signed(-32'she36b) : $signed(_GEN_3383); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3385 = 11'h538 == cnt[10:0] ? $signed(-32'she33c) : $signed(_GEN_3384); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3386 = 11'h539 == cnt[10:0] ? $signed(-32'she30e) : $signed(_GEN_3385); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3387 = 11'h53a == cnt[10:0] ? $signed(-32'she2df) : $signed(_GEN_3386); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3388 = 11'h53b == cnt[10:0] ? $signed(-32'she2b1) : $signed(_GEN_3387); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3389 = 11'h53c == cnt[10:0] ? $signed(-32'she282) : $signed(_GEN_3388); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3390 = 11'h53d == cnt[10:0] ? $signed(-32'she253) : $signed(_GEN_3389); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3391 = 11'h53e == cnt[10:0] ? $signed(-32'she224) : $signed(_GEN_3390); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3392 = 11'h53f == cnt[10:0] ? $signed(-32'she1f5) : $signed(_GEN_3391); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3393 = 11'h540 == cnt[10:0] ? $signed(-32'she1c6) : $signed(_GEN_3392); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3394 = 11'h541 == cnt[10:0] ? $signed(-32'she196) : $signed(_GEN_3393); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3395 = 11'h542 == cnt[10:0] ? $signed(-32'she167) : $signed(_GEN_3394); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3396 = 11'h543 == cnt[10:0] ? $signed(-32'she137) : $signed(_GEN_3395); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3397 = 11'h544 == cnt[10:0] ? $signed(-32'she107) : $signed(_GEN_3396); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3398 = 11'h545 == cnt[10:0] ? $signed(-32'she0d7) : $signed(_GEN_3397); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3399 = 11'h546 == cnt[10:0] ? $signed(-32'she0a7) : $signed(_GEN_3398); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3400 = 11'h547 == cnt[10:0] ? $signed(-32'she077) : $signed(_GEN_3399); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3401 = 11'h548 == cnt[10:0] ? $signed(-32'she046) : $signed(_GEN_3400); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3402 = 11'h549 == cnt[10:0] ? $signed(-32'she016) : $signed(_GEN_3401); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3403 = 11'h54a == cnt[10:0] ? $signed(-32'shdfe5) : $signed(_GEN_3402); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3404 = 11'h54b == cnt[10:0] ? $signed(-32'shdfb4) : $signed(_GEN_3403); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3405 = 11'h54c == cnt[10:0] ? $signed(-32'shdf83) : $signed(_GEN_3404); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3406 = 11'h54d == cnt[10:0] ? $signed(-32'shdf52) : $signed(_GEN_3405); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3407 = 11'h54e == cnt[10:0] ? $signed(-32'shdf21) : $signed(_GEN_3406); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3408 = 11'h54f == cnt[10:0] ? $signed(-32'shdef0) : $signed(_GEN_3407); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3409 = 11'h550 == cnt[10:0] ? $signed(-32'shdebe) : $signed(_GEN_3408); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3410 = 11'h551 == cnt[10:0] ? $signed(-32'shde8c) : $signed(_GEN_3409); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3411 = 11'h552 == cnt[10:0] ? $signed(-32'shde5b) : $signed(_GEN_3410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3412 = 11'h553 == cnt[10:0] ? $signed(-32'shde29) : $signed(_GEN_3411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3413 = 11'h554 == cnt[10:0] ? $signed(-32'shddf7) : $signed(_GEN_3412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3414 = 11'h555 == cnt[10:0] ? $signed(-32'shddc5) : $signed(_GEN_3413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3415 = 11'h556 == cnt[10:0] ? $signed(-32'shdd92) : $signed(_GEN_3414); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3416 = 11'h557 == cnt[10:0] ? $signed(-32'shdd60) : $signed(_GEN_3415); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3417 = 11'h558 == cnt[10:0] ? $signed(-32'shdd2d) : $signed(_GEN_3416); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3418 = 11'h559 == cnt[10:0] ? $signed(-32'shdcfb) : $signed(_GEN_3417); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3419 = 11'h55a == cnt[10:0] ? $signed(-32'shdcc8) : $signed(_GEN_3418); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3420 = 11'h55b == cnt[10:0] ? $signed(-32'shdc95) : $signed(_GEN_3419); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3421 = 11'h55c == cnt[10:0] ? $signed(-32'shdc62) : $signed(_GEN_3420); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3422 = 11'h55d == cnt[10:0] ? $signed(-32'shdc2f) : $signed(_GEN_3421); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3423 = 11'h55e == cnt[10:0] ? $signed(-32'shdbfb) : $signed(_GEN_3422); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3424 = 11'h55f == cnt[10:0] ? $signed(-32'shdbc8) : $signed(_GEN_3423); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3425 = 11'h560 == cnt[10:0] ? $signed(-32'shdb94) : $signed(_GEN_3424); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3426 = 11'h561 == cnt[10:0] ? $signed(-32'shdb60) : $signed(_GEN_3425); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3427 = 11'h562 == cnt[10:0] ? $signed(-32'shdb2c) : $signed(_GEN_3426); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3428 = 11'h563 == cnt[10:0] ? $signed(-32'shdaf8) : $signed(_GEN_3427); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3429 = 11'h564 == cnt[10:0] ? $signed(-32'shdac4) : $signed(_GEN_3428); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3430 = 11'h565 == cnt[10:0] ? $signed(-32'shda90) : $signed(_GEN_3429); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3431 = 11'h566 == cnt[10:0] ? $signed(-32'shda5c) : $signed(_GEN_3430); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3432 = 11'h567 == cnt[10:0] ? $signed(-32'shda27) : $signed(_GEN_3431); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3433 = 11'h568 == cnt[10:0] ? $signed(-32'shd9f2) : $signed(_GEN_3432); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3434 = 11'h569 == cnt[10:0] ? $signed(-32'shd9be) : $signed(_GEN_3433); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3435 = 11'h56a == cnt[10:0] ? $signed(-32'shd989) : $signed(_GEN_3434); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3436 = 11'h56b == cnt[10:0] ? $signed(-32'shd954) : $signed(_GEN_3435); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3437 = 11'h56c == cnt[10:0] ? $signed(-32'shd91e) : $signed(_GEN_3436); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3438 = 11'h56d == cnt[10:0] ? $signed(-32'shd8e9) : $signed(_GEN_3437); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3439 = 11'h56e == cnt[10:0] ? $signed(-32'shd8b4) : $signed(_GEN_3438); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3440 = 11'h56f == cnt[10:0] ? $signed(-32'shd87e) : $signed(_GEN_3439); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3441 = 11'h570 == cnt[10:0] ? $signed(-32'shd848) : $signed(_GEN_3440); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3442 = 11'h571 == cnt[10:0] ? $signed(-32'shd812) : $signed(_GEN_3441); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3443 = 11'h572 == cnt[10:0] ? $signed(-32'shd7dc) : $signed(_GEN_3442); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3444 = 11'h573 == cnt[10:0] ? $signed(-32'shd7a6) : $signed(_GEN_3443); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3445 = 11'h574 == cnt[10:0] ? $signed(-32'shd770) : $signed(_GEN_3444); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3446 = 11'h575 == cnt[10:0] ? $signed(-32'shd73a) : $signed(_GEN_3445); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3447 = 11'h576 == cnt[10:0] ? $signed(-32'shd703) : $signed(_GEN_3446); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3448 = 11'h577 == cnt[10:0] ? $signed(-32'shd6cd) : $signed(_GEN_3447); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3449 = 11'h578 == cnt[10:0] ? $signed(-32'shd696) : $signed(_GEN_3448); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3450 = 11'h579 == cnt[10:0] ? $signed(-32'shd65f) : $signed(_GEN_3449); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3451 = 11'h57a == cnt[10:0] ? $signed(-32'shd628) : $signed(_GEN_3450); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3452 = 11'h57b == cnt[10:0] ? $signed(-32'shd5f1) : $signed(_GEN_3451); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3453 = 11'h57c == cnt[10:0] ? $signed(-32'shd5ba) : $signed(_GEN_3452); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3454 = 11'h57d == cnt[10:0] ? $signed(-32'shd582) : $signed(_GEN_3453); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3455 = 11'h57e == cnt[10:0] ? $signed(-32'shd54b) : $signed(_GEN_3454); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3456 = 11'h57f == cnt[10:0] ? $signed(-32'shd513) : $signed(_GEN_3455); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3457 = 11'h580 == cnt[10:0] ? $signed(-32'shd4db) : $signed(_GEN_3456); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3458 = 11'h581 == cnt[10:0] ? $signed(-32'shd4a3) : $signed(_GEN_3457); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3459 = 11'h582 == cnt[10:0] ? $signed(-32'shd46b) : $signed(_GEN_3458); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3460 = 11'h583 == cnt[10:0] ? $signed(-32'shd433) : $signed(_GEN_3459); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3461 = 11'h584 == cnt[10:0] ? $signed(-32'shd3fb) : $signed(_GEN_3460); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3462 = 11'h585 == cnt[10:0] ? $signed(-32'shd3c2) : $signed(_GEN_3461); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3463 = 11'h586 == cnt[10:0] ? $signed(-32'shd38a) : $signed(_GEN_3462); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3464 = 11'h587 == cnt[10:0] ? $signed(-32'shd351) : $signed(_GEN_3463); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3465 = 11'h588 == cnt[10:0] ? $signed(-32'shd318) : $signed(_GEN_3464); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3466 = 11'h589 == cnt[10:0] ? $signed(-32'shd2df) : $signed(_GEN_3465); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3467 = 11'h58a == cnt[10:0] ? $signed(-32'shd2a6) : $signed(_GEN_3466); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3468 = 11'h58b == cnt[10:0] ? $signed(-32'shd26d) : $signed(_GEN_3467); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3469 = 11'h58c == cnt[10:0] ? $signed(-32'shd234) : $signed(_GEN_3468); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3470 = 11'h58d == cnt[10:0] ? $signed(-32'shd1fa) : $signed(_GEN_3469); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3471 = 11'h58e == cnt[10:0] ? $signed(-32'shd1c1) : $signed(_GEN_3470); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3472 = 11'h58f == cnt[10:0] ? $signed(-32'shd187) : $signed(_GEN_3471); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3473 = 11'h590 == cnt[10:0] ? $signed(-32'shd14d) : $signed(_GEN_3472); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3474 = 11'h591 == cnt[10:0] ? $signed(-32'shd113) : $signed(_GEN_3473); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3475 = 11'h592 == cnt[10:0] ? $signed(-32'shd0d9) : $signed(_GEN_3474); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3476 = 11'h593 == cnt[10:0] ? $signed(-32'shd09f) : $signed(_GEN_3475); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3477 = 11'h594 == cnt[10:0] ? $signed(-32'shd065) : $signed(_GEN_3476); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3478 = 11'h595 == cnt[10:0] ? $signed(-32'shd02a) : $signed(_GEN_3477); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3479 = 11'h596 == cnt[10:0] ? $signed(-32'shcff0) : $signed(_GEN_3478); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3480 = 11'h597 == cnt[10:0] ? $signed(-32'shcfb5) : $signed(_GEN_3479); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3481 = 11'h598 == cnt[10:0] ? $signed(-32'shcf7a) : $signed(_GEN_3480); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3482 = 11'h599 == cnt[10:0] ? $signed(-32'shcf3f) : $signed(_GEN_3481); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3483 = 11'h59a == cnt[10:0] ? $signed(-32'shcf04) : $signed(_GEN_3482); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3484 = 11'h59b == cnt[10:0] ? $signed(-32'shcec9) : $signed(_GEN_3483); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3485 = 11'h59c == cnt[10:0] ? $signed(-32'shce8e) : $signed(_GEN_3484); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3486 = 11'h59d == cnt[10:0] ? $signed(-32'shce52) : $signed(_GEN_3485); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3487 = 11'h59e == cnt[10:0] ? $signed(-32'shce17) : $signed(_GEN_3486); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3488 = 11'h59f == cnt[10:0] ? $signed(-32'shcddb) : $signed(_GEN_3487); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3489 = 11'h5a0 == cnt[10:0] ? $signed(-32'shcd9f) : $signed(_GEN_3488); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3490 = 11'h5a1 == cnt[10:0] ? $signed(-32'shcd63) : $signed(_GEN_3489); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3491 = 11'h5a2 == cnt[10:0] ? $signed(-32'shcd27) : $signed(_GEN_3490); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3492 = 11'h5a3 == cnt[10:0] ? $signed(-32'shcceb) : $signed(_GEN_3491); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3493 = 11'h5a4 == cnt[10:0] ? $signed(-32'shccae) : $signed(_GEN_3492); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3494 = 11'h5a5 == cnt[10:0] ? $signed(-32'shcc72) : $signed(_GEN_3493); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3495 = 11'h5a6 == cnt[10:0] ? $signed(-32'shcc35) : $signed(_GEN_3494); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3496 = 11'h5a7 == cnt[10:0] ? $signed(-32'shcbf9) : $signed(_GEN_3495); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3497 = 11'h5a8 == cnt[10:0] ? $signed(-32'shcbbc) : $signed(_GEN_3496); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3498 = 11'h5a9 == cnt[10:0] ? $signed(-32'shcb7f) : $signed(_GEN_3497); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3499 = 11'h5aa == cnt[10:0] ? $signed(-32'shcb42) : $signed(_GEN_3498); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3500 = 11'h5ab == cnt[10:0] ? $signed(-32'shcb05) : $signed(_GEN_3499); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3501 = 11'h5ac == cnt[10:0] ? $signed(-32'shcac7) : $signed(_GEN_3500); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3502 = 11'h5ad == cnt[10:0] ? $signed(-32'shca8a) : $signed(_GEN_3501); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3503 = 11'h5ae == cnt[10:0] ? $signed(-32'shca4d) : $signed(_GEN_3502); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3504 = 11'h5af == cnt[10:0] ? $signed(-32'shca0f) : $signed(_GEN_3503); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3505 = 11'h5b0 == cnt[10:0] ? $signed(-32'shc9d1) : $signed(_GEN_3504); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3506 = 11'h5b1 == cnt[10:0] ? $signed(-32'shc993) : $signed(_GEN_3505); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3507 = 11'h5b2 == cnt[10:0] ? $signed(-32'shc955) : $signed(_GEN_3506); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3508 = 11'h5b3 == cnt[10:0] ? $signed(-32'shc917) : $signed(_GEN_3507); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3509 = 11'h5b4 == cnt[10:0] ? $signed(-32'shc8d9) : $signed(_GEN_3508); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3510 = 11'h5b5 == cnt[10:0] ? $signed(-32'shc89a) : $signed(_GEN_3509); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3511 = 11'h5b6 == cnt[10:0] ? $signed(-32'shc85c) : $signed(_GEN_3510); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3512 = 11'h5b7 == cnt[10:0] ? $signed(-32'shc81d) : $signed(_GEN_3511); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3513 = 11'h5b8 == cnt[10:0] ? $signed(-32'shc7de) : $signed(_GEN_3512); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3514 = 11'h5b9 == cnt[10:0] ? $signed(-32'shc7a0) : $signed(_GEN_3513); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3515 = 11'h5ba == cnt[10:0] ? $signed(-32'shc761) : $signed(_GEN_3514); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3516 = 11'h5bb == cnt[10:0] ? $signed(-32'shc721) : $signed(_GEN_3515); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3517 = 11'h5bc == cnt[10:0] ? $signed(-32'shc6e2) : $signed(_GEN_3516); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3518 = 11'h5bd == cnt[10:0] ? $signed(-32'shc6a3) : $signed(_GEN_3517); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3519 = 11'h5be == cnt[10:0] ? $signed(-32'shc663) : $signed(_GEN_3518); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3520 = 11'h5bf == cnt[10:0] ? $signed(-32'shc624) : $signed(_GEN_3519); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3521 = 11'h5c0 == cnt[10:0] ? $signed(-32'shc5e4) : $signed(_GEN_3520); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3522 = 11'h5c1 == cnt[10:0] ? $signed(-32'shc5a4) : $signed(_GEN_3521); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3523 = 11'h5c2 == cnt[10:0] ? $signed(-32'shc564) : $signed(_GEN_3522); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3524 = 11'h5c3 == cnt[10:0] ? $signed(-32'shc524) : $signed(_GEN_3523); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3525 = 11'h5c4 == cnt[10:0] ? $signed(-32'shc4e4) : $signed(_GEN_3524); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3526 = 11'h5c5 == cnt[10:0] ? $signed(-32'shc4a4) : $signed(_GEN_3525); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3527 = 11'h5c6 == cnt[10:0] ? $signed(-32'shc463) : $signed(_GEN_3526); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3528 = 11'h5c7 == cnt[10:0] ? $signed(-32'shc423) : $signed(_GEN_3527); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3529 = 11'h5c8 == cnt[10:0] ? $signed(-32'shc3e2) : $signed(_GEN_3528); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3530 = 11'h5c9 == cnt[10:0] ? $signed(-32'shc3a1) : $signed(_GEN_3529); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3531 = 11'h5ca == cnt[10:0] ? $signed(-32'shc360) : $signed(_GEN_3530); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3532 = 11'h5cb == cnt[10:0] ? $signed(-32'shc31f) : $signed(_GEN_3531); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3533 = 11'h5cc == cnt[10:0] ? $signed(-32'shc2de) : $signed(_GEN_3532); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3534 = 11'h5cd == cnt[10:0] ? $signed(-32'shc29d) : $signed(_GEN_3533); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3535 = 11'h5ce == cnt[10:0] ? $signed(-32'shc25c) : $signed(_GEN_3534); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3536 = 11'h5cf == cnt[10:0] ? $signed(-32'shc21a) : $signed(_GEN_3535); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3537 = 11'h5d0 == cnt[10:0] ? $signed(-32'shc1d8) : $signed(_GEN_3536); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3538 = 11'h5d1 == cnt[10:0] ? $signed(-32'shc197) : $signed(_GEN_3537); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3539 = 11'h5d2 == cnt[10:0] ? $signed(-32'shc155) : $signed(_GEN_3538); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3540 = 11'h5d3 == cnt[10:0] ? $signed(-32'shc113) : $signed(_GEN_3539); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3541 = 11'h5d4 == cnt[10:0] ? $signed(-32'shc0d1) : $signed(_GEN_3540); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3542 = 11'h5d5 == cnt[10:0] ? $signed(-32'shc08f) : $signed(_GEN_3541); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3543 = 11'h5d6 == cnt[10:0] ? $signed(-32'shc04c) : $signed(_GEN_3542); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3544 = 11'h5d7 == cnt[10:0] ? $signed(-32'shc00a) : $signed(_GEN_3543); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3545 = 11'h5d8 == cnt[10:0] ? $signed(-32'shbfc7) : $signed(_GEN_3544); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3546 = 11'h5d9 == cnt[10:0] ? $signed(-32'shbf85) : $signed(_GEN_3545); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3547 = 11'h5da == cnt[10:0] ? $signed(-32'shbf42) : $signed(_GEN_3546); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3548 = 11'h5db == cnt[10:0] ? $signed(-32'shbeff) : $signed(_GEN_3547); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3549 = 11'h5dc == cnt[10:0] ? $signed(-32'shbebc) : $signed(_GEN_3548); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3550 = 11'h5dd == cnt[10:0] ? $signed(-32'shbe79) : $signed(_GEN_3549); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3551 = 11'h5de == cnt[10:0] ? $signed(-32'shbe36) : $signed(_GEN_3550); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3552 = 11'h5df == cnt[10:0] ? $signed(-32'shbdf2) : $signed(_GEN_3551); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3553 = 11'h5e0 == cnt[10:0] ? $signed(-32'shbdaf) : $signed(_GEN_3552); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3554 = 11'h5e1 == cnt[10:0] ? $signed(-32'shbd6b) : $signed(_GEN_3553); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3555 = 11'h5e2 == cnt[10:0] ? $signed(-32'shbd28) : $signed(_GEN_3554); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3556 = 11'h5e3 == cnt[10:0] ? $signed(-32'shbce4) : $signed(_GEN_3555); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3557 = 11'h5e4 == cnt[10:0] ? $signed(-32'shbca0) : $signed(_GEN_3556); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3558 = 11'h5e5 == cnt[10:0] ? $signed(-32'shbc5c) : $signed(_GEN_3557); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3559 = 11'h5e6 == cnt[10:0] ? $signed(-32'shbc18) : $signed(_GEN_3558); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3560 = 11'h5e7 == cnt[10:0] ? $signed(-32'shbbd4) : $signed(_GEN_3559); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3561 = 11'h5e8 == cnt[10:0] ? $signed(-32'shbb8f) : $signed(_GEN_3560); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3562 = 11'h5e9 == cnt[10:0] ? $signed(-32'shbb4b) : $signed(_GEN_3561); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3563 = 11'h5ea == cnt[10:0] ? $signed(-32'shbb06) : $signed(_GEN_3562); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3564 = 11'h5eb == cnt[10:0] ? $signed(-32'shbac1) : $signed(_GEN_3563); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3565 = 11'h5ec == cnt[10:0] ? $signed(-32'shba7d) : $signed(_GEN_3564); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3566 = 11'h5ed == cnt[10:0] ? $signed(-32'shba38) : $signed(_GEN_3565); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3567 = 11'h5ee == cnt[10:0] ? $signed(-32'shb9f3) : $signed(_GEN_3566); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3568 = 11'h5ef == cnt[10:0] ? $signed(-32'shb9ae) : $signed(_GEN_3567); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3569 = 11'h5f0 == cnt[10:0] ? $signed(-32'shb968) : $signed(_GEN_3568); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3570 = 11'h5f1 == cnt[10:0] ? $signed(-32'shb923) : $signed(_GEN_3569); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3571 = 11'h5f2 == cnt[10:0] ? $signed(-32'shb8dd) : $signed(_GEN_3570); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3572 = 11'h5f3 == cnt[10:0] ? $signed(-32'shb898) : $signed(_GEN_3571); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3573 = 11'h5f4 == cnt[10:0] ? $signed(-32'shb852) : $signed(_GEN_3572); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3574 = 11'h5f5 == cnt[10:0] ? $signed(-32'shb80c) : $signed(_GEN_3573); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3575 = 11'h5f6 == cnt[10:0] ? $signed(-32'shb7c6) : $signed(_GEN_3574); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3576 = 11'h5f7 == cnt[10:0] ? $signed(-32'shb780) : $signed(_GEN_3575); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3577 = 11'h5f8 == cnt[10:0] ? $signed(-32'shb73a) : $signed(_GEN_3576); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3578 = 11'h5f9 == cnt[10:0] ? $signed(-32'shb6f4) : $signed(_GEN_3577); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3579 = 11'h5fa == cnt[10:0] ? $signed(-32'shb6ad) : $signed(_GEN_3578); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3580 = 11'h5fb == cnt[10:0] ? $signed(-32'shb667) : $signed(_GEN_3579); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3581 = 11'h5fc == cnt[10:0] ? $signed(-32'shb620) : $signed(_GEN_3580); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3582 = 11'h5fd == cnt[10:0] ? $signed(-32'shb5da) : $signed(_GEN_3581); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3583 = 11'h5fe == cnt[10:0] ? $signed(-32'shb593) : $signed(_GEN_3582); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3584 = 11'h5ff == cnt[10:0] ? $signed(-32'shb54c) : $signed(_GEN_3583); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3585 = 11'h600 == cnt[10:0] ? $signed(-32'shb505) : $signed(_GEN_3584); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3586 = 11'h601 == cnt[10:0] ? $signed(-32'shb4be) : $signed(_GEN_3585); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3587 = 11'h602 == cnt[10:0] ? $signed(-32'shb477) : $signed(_GEN_3586); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3588 = 11'h603 == cnt[10:0] ? $signed(-32'shb42f) : $signed(_GEN_3587); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3589 = 11'h604 == cnt[10:0] ? $signed(-32'shb3e8) : $signed(_GEN_3588); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3590 = 11'h605 == cnt[10:0] ? $signed(-32'shb3a0) : $signed(_GEN_3589); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3591 = 11'h606 == cnt[10:0] ? $signed(-32'shb358) : $signed(_GEN_3590); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3592 = 11'h607 == cnt[10:0] ? $signed(-32'shb311) : $signed(_GEN_3591); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3593 = 11'h608 == cnt[10:0] ? $signed(-32'shb2c9) : $signed(_GEN_3592); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3594 = 11'h609 == cnt[10:0] ? $signed(-32'shb281) : $signed(_GEN_3593); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3595 = 11'h60a == cnt[10:0] ? $signed(-32'shb239) : $signed(_GEN_3594); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3596 = 11'h60b == cnt[10:0] ? $signed(-32'shb1f0) : $signed(_GEN_3595); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3597 = 11'h60c == cnt[10:0] ? $signed(-32'shb1a8) : $signed(_GEN_3596); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3598 = 11'h60d == cnt[10:0] ? $signed(-32'shb160) : $signed(_GEN_3597); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3599 = 11'h60e == cnt[10:0] ? $signed(-32'shb117) : $signed(_GEN_3598); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3600 = 11'h60f == cnt[10:0] ? $signed(-32'shb0ce) : $signed(_GEN_3599); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3601 = 11'h610 == cnt[10:0] ? $signed(-32'shb086) : $signed(_GEN_3600); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3602 = 11'h611 == cnt[10:0] ? $signed(-32'shb03d) : $signed(_GEN_3601); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3603 = 11'h612 == cnt[10:0] ? $signed(-32'shaff4) : $signed(_GEN_3602); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3604 = 11'h613 == cnt[10:0] ? $signed(-32'shafab) : $signed(_GEN_3603); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3605 = 11'h614 == cnt[10:0] ? $signed(-32'shaf62) : $signed(_GEN_3604); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3606 = 11'h615 == cnt[10:0] ? $signed(-32'shaf18) : $signed(_GEN_3605); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3607 = 11'h616 == cnt[10:0] ? $signed(-32'shaecf) : $signed(_GEN_3606); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3608 = 11'h617 == cnt[10:0] ? $signed(-32'shae85) : $signed(_GEN_3607); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3609 = 11'h618 == cnt[10:0] ? $signed(-32'shae3c) : $signed(_GEN_3608); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3610 = 11'h619 == cnt[10:0] ? $signed(-32'shadf2) : $signed(_GEN_3609); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3611 = 11'h61a == cnt[10:0] ? $signed(-32'shada8) : $signed(_GEN_3610); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3612 = 11'h61b == cnt[10:0] ? $signed(-32'shad5e) : $signed(_GEN_3611); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3613 = 11'h61c == cnt[10:0] ? $signed(-32'shad14) : $signed(_GEN_3612); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3614 = 11'h61d == cnt[10:0] ? $signed(-32'shacca) : $signed(_GEN_3613); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3615 = 11'h61e == cnt[10:0] ? $signed(-32'shac80) : $signed(_GEN_3614); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3616 = 11'h61f == cnt[10:0] ? $signed(-32'shac36) : $signed(_GEN_3615); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3617 = 11'h620 == cnt[10:0] ? $signed(-32'shabeb) : $signed(_GEN_3616); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3618 = 11'h621 == cnt[10:0] ? $signed(-32'shaba1) : $signed(_GEN_3617); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3619 = 11'h622 == cnt[10:0] ? $signed(-32'shab56) : $signed(_GEN_3618); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3620 = 11'h623 == cnt[10:0] ? $signed(-32'shab0b) : $signed(_GEN_3619); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3621 = 11'h624 == cnt[10:0] ? $signed(-32'shaac1) : $signed(_GEN_3620); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3622 = 11'h625 == cnt[10:0] ? $signed(-32'shaa76) : $signed(_GEN_3621); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3623 = 11'h626 == cnt[10:0] ? $signed(-32'shaa2a) : $signed(_GEN_3622); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3624 = 11'h627 == cnt[10:0] ? $signed(-32'sha9df) : $signed(_GEN_3623); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3625 = 11'h628 == cnt[10:0] ? $signed(-32'sha994) : $signed(_GEN_3624); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3626 = 11'h629 == cnt[10:0] ? $signed(-32'sha949) : $signed(_GEN_3625); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3627 = 11'h62a == cnt[10:0] ? $signed(-32'sha8fd) : $signed(_GEN_3626); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3628 = 11'h62b == cnt[10:0] ? $signed(-32'sha8b2) : $signed(_GEN_3627); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3629 = 11'h62c == cnt[10:0] ? $signed(-32'sha866) : $signed(_GEN_3628); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3630 = 11'h62d == cnt[10:0] ? $signed(-32'sha81a) : $signed(_GEN_3629); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3631 = 11'h62e == cnt[10:0] ? $signed(-32'sha7ce) : $signed(_GEN_3630); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3632 = 11'h62f == cnt[10:0] ? $signed(-32'sha782) : $signed(_GEN_3631); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3633 = 11'h630 == cnt[10:0] ? $signed(-32'sha736) : $signed(_GEN_3632); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3634 = 11'h631 == cnt[10:0] ? $signed(-32'sha6ea) : $signed(_GEN_3633); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3635 = 11'h632 == cnt[10:0] ? $signed(-32'sha69e) : $signed(_GEN_3634); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3636 = 11'h633 == cnt[10:0] ? $signed(-32'sha652) : $signed(_GEN_3635); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3637 = 11'h634 == cnt[10:0] ? $signed(-32'sha605) : $signed(_GEN_3636); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3638 = 11'h635 == cnt[10:0] ? $signed(-32'sha5b8) : $signed(_GEN_3637); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3639 = 11'h636 == cnt[10:0] ? $signed(-32'sha56c) : $signed(_GEN_3638); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3640 = 11'h637 == cnt[10:0] ? $signed(-32'sha51f) : $signed(_GEN_3639); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3641 = 11'h638 == cnt[10:0] ? $signed(-32'sha4d2) : $signed(_GEN_3640); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3642 = 11'h639 == cnt[10:0] ? $signed(-32'sha485) : $signed(_GEN_3641); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3643 = 11'h63a == cnt[10:0] ? $signed(-32'sha438) : $signed(_GEN_3642); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3644 = 11'h63b == cnt[10:0] ? $signed(-32'sha3eb) : $signed(_GEN_3643); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3645 = 11'h63c == cnt[10:0] ? $signed(-32'sha39e) : $signed(_GEN_3644); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3646 = 11'h63d == cnt[10:0] ? $signed(-32'sha350) : $signed(_GEN_3645); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3647 = 11'h63e == cnt[10:0] ? $signed(-32'sha303) : $signed(_GEN_3646); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3648 = 11'h63f == cnt[10:0] ? $signed(-32'sha2b5) : $signed(_GEN_3647); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3649 = 11'h640 == cnt[10:0] ? $signed(-32'sha268) : $signed(_GEN_3648); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3650 = 11'h641 == cnt[10:0] ? $signed(-32'sha21a) : $signed(_GEN_3649); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3651 = 11'h642 == cnt[10:0] ? $signed(-32'sha1cc) : $signed(_GEN_3650); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3652 = 11'h643 == cnt[10:0] ? $signed(-32'sha17e) : $signed(_GEN_3651); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3653 = 11'h644 == cnt[10:0] ? $signed(-32'sha130) : $signed(_GEN_3652); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3654 = 11'h645 == cnt[10:0] ? $signed(-32'sha0e2) : $signed(_GEN_3653); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3655 = 11'h646 == cnt[10:0] ? $signed(-32'sha094) : $signed(_GEN_3654); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3656 = 11'h647 == cnt[10:0] ? $signed(-32'sha045) : $signed(_GEN_3655); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3657 = 11'h648 == cnt[10:0] ? $signed(-32'sh9ff7) : $signed(_GEN_3656); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3658 = 11'h649 == cnt[10:0] ? $signed(-32'sh9fa8) : $signed(_GEN_3657); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3659 = 11'h64a == cnt[10:0] ? $signed(-32'sh9f5a) : $signed(_GEN_3658); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3660 = 11'h64b == cnt[10:0] ? $signed(-32'sh9f0b) : $signed(_GEN_3659); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3661 = 11'h64c == cnt[10:0] ? $signed(-32'sh9ebc) : $signed(_GEN_3660); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3662 = 11'h64d == cnt[10:0] ? $signed(-32'sh9e6d) : $signed(_GEN_3661); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3663 = 11'h64e == cnt[10:0] ? $signed(-32'sh9e1e) : $signed(_GEN_3662); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3664 = 11'h64f == cnt[10:0] ? $signed(-32'sh9dcf) : $signed(_GEN_3663); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3665 = 11'h650 == cnt[10:0] ? $signed(-32'sh9d80) : $signed(_GEN_3664); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3666 = 11'h651 == cnt[10:0] ? $signed(-32'sh9d31) : $signed(_GEN_3665); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3667 = 11'h652 == cnt[10:0] ? $signed(-32'sh9ce1) : $signed(_GEN_3666); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3668 = 11'h653 == cnt[10:0] ? $signed(-32'sh9c92) : $signed(_GEN_3667); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3669 = 11'h654 == cnt[10:0] ? $signed(-32'sh9c42) : $signed(_GEN_3668); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3670 = 11'h655 == cnt[10:0] ? $signed(-32'sh9bf2) : $signed(_GEN_3669); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3671 = 11'h656 == cnt[10:0] ? $signed(-32'sh9ba3) : $signed(_GEN_3670); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3672 = 11'h657 == cnt[10:0] ? $signed(-32'sh9b53) : $signed(_GEN_3671); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3673 = 11'h658 == cnt[10:0] ? $signed(-32'sh9b03) : $signed(_GEN_3672); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3674 = 11'h659 == cnt[10:0] ? $signed(-32'sh9ab3) : $signed(_GEN_3673); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3675 = 11'h65a == cnt[10:0] ? $signed(-32'sh9a63) : $signed(_GEN_3674); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3676 = 11'h65b == cnt[10:0] ? $signed(-32'sh9a12) : $signed(_GEN_3675); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3677 = 11'h65c == cnt[10:0] ? $signed(-32'sh99c2) : $signed(_GEN_3676); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3678 = 11'h65d == cnt[10:0] ? $signed(-32'sh9972) : $signed(_GEN_3677); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3679 = 11'h65e == cnt[10:0] ? $signed(-32'sh9921) : $signed(_GEN_3678); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3680 = 11'h65f == cnt[10:0] ? $signed(-32'sh98d0) : $signed(_GEN_3679); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3681 = 11'h660 == cnt[10:0] ? $signed(-32'sh9880) : $signed(_GEN_3680); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3682 = 11'h661 == cnt[10:0] ? $signed(-32'sh982f) : $signed(_GEN_3681); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3683 = 11'h662 == cnt[10:0] ? $signed(-32'sh97de) : $signed(_GEN_3682); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3684 = 11'h663 == cnt[10:0] ? $signed(-32'sh978d) : $signed(_GEN_3683); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3685 = 11'h664 == cnt[10:0] ? $signed(-32'sh973c) : $signed(_GEN_3684); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3686 = 11'h665 == cnt[10:0] ? $signed(-32'sh96eb) : $signed(_GEN_3685); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3687 = 11'h666 == cnt[10:0] ? $signed(-32'sh969a) : $signed(_GEN_3686); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3688 = 11'h667 == cnt[10:0] ? $signed(-32'sh9648) : $signed(_GEN_3687); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3689 = 11'h668 == cnt[10:0] ? $signed(-32'sh95f7) : $signed(_GEN_3688); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3690 = 11'h669 == cnt[10:0] ? $signed(-32'sh95a5) : $signed(_GEN_3689); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3691 = 11'h66a == cnt[10:0] ? $signed(-32'sh9554) : $signed(_GEN_3690); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3692 = 11'h66b == cnt[10:0] ? $signed(-32'sh9502) : $signed(_GEN_3691); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3693 = 11'h66c == cnt[10:0] ? $signed(-32'sh94b0) : $signed(_GEN_3692); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3694 = 11'h66d == cnt[10:0] ? $signed(-32'sh945e) : $signed(_GEN_3693); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3695 = 11'h66e == cnt[10:0] ? $signed(-32'sh940c) : $signed(_GEN_3694); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3696 = 11'h66f == cnt[10:0] ? $signed(-32'sh93ba) : $signed(_GEN_3695); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3697 = 11'h670 == cnt[10:0] ? $signed(-32'sh9368) : $signed(_GEN_3696); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3698 = 11'h671 == cnt[10:0] ? $signed(-32'sh9316) : $signed(_GEN_3697); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3699 = 11'h672 == cnt[10:0] ? $signed(-32'sh92c4) : $signed(_GEN_3698); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3700 = 11'h673 == cnt[10:0] ? $signed(-32'sh9271) : $signed(_GEN_3699); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3701 = 11'h674 == cnt[10:0] ? $signed(-32'sh921f) : $signed(_GEN_3700); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3702 = 11'h675 == cnt[10:0] ? $signed(-32'sh91cc) : $signed(_GEN_3701); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3703 = 11'h676 == cnt[10:0] ? $signed(-32'sh9179) : $signed(_GEN_3702); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3704 = 11'h677 == cnt[10:0] ? $signed(-32'sh9127) : $signed(_GEN_3703); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3705 = 11'h678 == cnt[10:0] ? $signed(-32'sh90d4) : $signed(_GEN_3704); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3706 = 11'h679 == cnt[10:0] ? $signed(-32'sh9081) : $signed(_GEN_3705); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3707 = 11'h67a == cnt[10:0] ? $signed(-32'sh902e) : $signed(_GEN_3706); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3708 = 11'h67b == cnt[10:0] ? $signed(-32'sh8fdb) : $signed(_GEN_3707); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3709 = 11'h67c == cnt[10:0] ? $signed(-32'sh8f88) : $signed(_GEN_3708); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3710 = 11'h67d == cnt[10:0] ? $signed(-32'sh8f34) : $signed(_GEN_3709); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3711 = 11'h67e == cnt[10:0] ? $signed(-32'sh8ee1) : $signed(_GEN_3710); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3712 = 11'h67f == cnt[10:0] ? $signed(-32'sh8e8d) : $signed(_GEN_3711); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3713 = 11'h680 == cnt[10:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3712); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3714 = 11'h681 == cnt[10:0] ? $signed(-32'sh8de6) : $signed(_GEN_3713); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3715 = 11'h682 == cnt[10:0] ? $signed(-32'sh8d93) : $signed(_GEN_3714); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3716 = 11'h683 == cnt[10:0] ? $signed(-32'sh8d3f) : $signed(_GEN_3715); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3717 = 11'h684 == cnt[10:0] ? $signed(-32'sh8ceb) : $signed(_GEN_3716); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3718 = 11'h685 == cnt[10:0] ? $signed(-32'sh8c97) : $signed(_GEN_3717); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3719 = 11'h686 == cnt[10:0] ? $signed(-32'sh8c43) : $signed(_GEN_3718); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3720 = 11'h687 == cnt[10:0] ? $signed(-32'sh8bef) : $signed(_GEN_3719); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3721 = 11'h688 == cnt[10:0] ? $signed(-32'sh8b9a) : $signed(_GEN_3720); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3722 = 11'h689 == cnt[10:0] ? $signed(-32'sh8b46) : $signed(_GEN_3721); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3723 = 11'h68a == cnt[10:0] ? $signed(-32'sh8af2) : $signed(_GEN_3722); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3724 = 11'h68b == cnt[10:0] ? $signed(-32'sh8a9d) : $signed(_GEN_3723); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3725 = 11'h68c == cnt[10:0] ? $signed(-32'sh8a49) : $signed(_GEN_3724); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3726 = 11'h68d == cnt[10:0] ? $signed(-32'sh89f4) : $signed(_GEN_3725); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3727 = 11'h68e == cnt[10:0] ? $signed(-32'sh899f) : $signed(_GEN_3726); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3728 = 11'h68f == cnt[10:0] ? $signed(-32'sh894a) : $signed(_GEN_3727); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3729 = 11'h690 == cnt[10:0] ? $signed(-32'sh88f6) : $signed(_GEN_3728); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3730 = 11'h691 == cnt[10:0] ? $signed(-32'sh88a1) : $signed(_GEN_3729); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3731 = 11'h692 == cnt[10:0] ? $signed(-32'sh884c) : $signed(_GEN_3730); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3732 = 11'h693 == cnt[10:0] ? $signed(-32'sh87f6) : $signed(_GEN_3731); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3733 = 11'h694 == cnt[10:0] ? $signed(-32'sh87a1) : $signed(_GEN_3732); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3734 = 11'h695 == cnt[10:0] ? $signed(-32'sh874c) : $signed(_GEN_3733); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3735 = 11'h696 == cnt[10:0] ? $signed(-32'sh86f7) : $signed(_GEN_3734); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3736 = 11'h697 == cnt[10:0] ? $signed(-32'sh86a1) : $signed(_GEN_3735); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3737 = 11'h698 == cnt[10:0] ? $signed(-32'sh864c) : $signed(_GEN_3736); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3738 = 11'h699 == cnt[10:0] ? $signed(-32'sh85f6) : $signed(_GEN_3737); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3739 = 11'h69a == cnt[10:0] ? $signed(-32'sh85a0) : $signed(_GEN_3738); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3740 = 11'h69b == cnt[10:0] ? $signed(-32'sh854a) : $signed(_GEN_3739); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3741 = 11'h69c == cnt[10:0] ? $signed(-32'sh84f5) : $signed(_GEN_3740); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3742 = 11'h69d == cnt[10:0] ? $signed(-32'sh849f) : $signed(_GEN_3741); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3743 = 11'h69e == cnt[10:0] ? $signed(-32'sh8449) : $signed(_GEN_3742); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3744 = 11'h69f == cnt[10:0] ? $signed(-32'sh83f2) : $signed(_GEN_3743); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3745 = 11'h6a0 == cnt[10:0] ? $signed(-32'sh839c) : $signed(_GEN_3744); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3746 = 11'h6a1 == cnt[10:0] ? $signed(-32'sh8346) : $signed(_GEN_3745); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3747 = 11'h6a2 == cnt[10:0] ? $signed(-32'sh82f0) : $signed(_GEN_3746); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3748 = 11'h6a3 == cnt[10:0] ? $signed(-32'sh8299) : $signed(_GEN_3747); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3749 = 11'h6a4 == cnt[10:0] ? $signed(-32'sh8243) : $signed(_GEN_3748); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3750 = 11'h6a5 == cnt[10:0] ? $signed(-32'sh81ec) : $signed(_GEN_3749); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3751 = 11'h6a6 == cnt[10:0] ? $signed(-32'sh8195) : $signed(_GEN_3750); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3752 = 11'h6a7 == cnt[10:0] ? $signed(-32'sh813f) : $signed(_GEN_3751); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3753 = 11'h6a8 == cnt[10:0] ? $signed(-32'sh80e8) : $signed(_GEN_3752); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3754 = 11'h6a9 == cnt[10:0] ? $signed(-32'sh8091) : $signed(_GEN_3753); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3755 = 11'h6aa == cnt[10:0] ? $signed(-32'sh803a) : $signed(_GEN_3754); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3756 = 11'h6ab == cnt[10:0] ? $signed(-32'sh7fe3) : $signed(_GEN_3755); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3757 = 11'h6ac == cnt[10:0] ? $signed(-32'sh7f8c) : $signed(_GEN_3756); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3758 = 11'h6ad == cnt[10:0] ? $signed(-32'sh7f35) : $signed(_GEN_3757); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3759 = 11'h6ae == cnt[10:0] ? $signed(-32'sh7edd) : $signed(_GEN_3758); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3760 = 11'h6af == cnt[10:0] ? $signed(-32'sh7e86) : $signed(_GEN_3759); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3761 = 11'h6b0 == cnt[10:0] ? $signed(-32'sh7e2f) : $signed(_GEN_3760); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3762 = 11'h6b1 == cnt[10:0] ? $signed(-32'sh7dd7) : $signed(_GEN_3761); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3763 = 11'h6b2 == cnt[10:0] ? $signed(-32'sh7d7f) : $signed(_GEN_3762); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3764 = 11'h6b3 == cnt[10:0] ? $signed(-32'sh7d28) : $signed(_GEN_3763); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3765 = 11'h6b4 == cnt[10:0] ? $signed(-32'sh7cd0) : $signed(_GEN_3764); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3766 = 11'h6b5 == cnt[10:0] ? $signed(-32'sh7c78) : $signed(_GEN_3765); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3767 = 11'h6b6 == cnt[10:0] ? $signed(-32'sh7c20) : $signed(_GEN_3766); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3768 = 11'h6b7 == cnt[10:0] ? $signed(-32'sh7bc8) : $signed(_GEN_3767); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3769 = 11'h6b8 == cnt[10:0] ? $signed(-32'sh7b70) : $signed(_GEN_3768); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3770 = 11'h6b9 == cnt[10:0] ? $signed(-32'sh7b18) : $signed(_GEN_3769); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3771 = 11'h6ba == cnt[10:0] ? $signed(-32'sh7ac0) : $signed(_GEN_3770); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3772 = 11'h6bb == cnt[10:0] ? $signed(-32'sh7a68) : $signed(_GEN_3771); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3773 = 11'h6bc == cnt[10:0] ? $signed(-32'sh7a10) : $signed(_GEN_3772); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3774 = 11'h6bd == cnt[10:0] ? $signed(-32'sh79b7) : $signed(_GEN_3773); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3775 = 11'h6be == cnt[10:0] ? $signed(-32'sh795f) : $signed(_GEN_3774); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3776 = 11'h6bf == cnt[10:0] ? $signed(-32'sh7906) : $signed(_GEN_3775); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3777 = 11'h6c0 == cnt[10:0] ? $signed(-32'sh78ad) : $signed(_GEN_3776); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3778 = 11'h6c1 == cnt[10:0] ? $signed(-32'sh7855) : $signed(_GEN_3777); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3779 = 11'h6c2 == cnt[10:0] ? $signed(-32'sh77fc) : $signed(_GEN_3778); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3780 = 11'h6c3 == cnt[10:0] ? $signed(-32'sh77a3) : $signed(_GEN_3779); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3781 = 11'h6c4 == cnt[10:0] ? $signed(-32'sh774a) : $signed(_GEN_3780); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3782 = 11'h6c5 == cnt[10:0] ? $signed(-32'sh76f1) : $signed(_GEN_3781); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3783 = 11'h6c6 == cnt[10:0] ? $signed(-32'sh7698) : $signed(_GEN_3782); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3784 = 11'h6c7 == cnt[10:0] ? $signed(-32'sh763f) : $signed(_GEN_3783); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3785 = 11'h6c8 == cnt[10:0] ? $signed(-32'sh75e6) : $signed(_GEN_3784); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3786 = 11'h6c9 == cnt[10:0] ? $signed(-32'sh758d) : $signed(_GEN_3785); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3787 = 11'h6ca == cnt[10:0] ? $signed(-32'sh7533) : $signed(_GEN_3786); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3788 = 11'h6cb == cnt[10:0] ? $signed(-32'sh74da) : $signed(_GEN_3787); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3789 = 11'h6cc == cnt[10:0] ? $signed(-32'sh7480) : $signed(_GEN_3788); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3790 = 11'h6cd == cnt[10:0] ? $signed(-32'sh7427) : $signed(_GEN_3789); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3791 = 11'h6ce == cnt[10:0] ? $signed(-32'sh73cd) : $signed(_GEN_3790); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3792 = 11'h6cf == cnt[10:0] ? $signed(-32'sh7373) : $signed(_GEN_3791); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3793 = 11'h6d0 == cnt[10:0] ? $signed(-32'sh731a) : $signed(_GEN_3792); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3794 = 11'h6d1 == cnt[10:0] ? $signed(-32'sh72c0) : $signed(_GEN_3793); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3795 = 11'h6d2 == cnt[10:0] ? $signed(-32'sh7266) : $signed(_GEN_3794); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3796 = 11'h6d3 == cnt[10:0] ? $signed(-32'sh720c) : $signed(_GEN_3795); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3797 = 11'h6d4 == cnt[10:0] ? $signed(-32'sh71b2) : $signed(_GEN_3796); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3798 = 11'h6d5 == cnt[10:0] ? $signed(-32'sh7158) : $signed(_GEN_3797); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3799 = 11'h6d6 == cnt[10:0] ? $signed(-32'sh70fe) : $signed(_GEN_3798); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3800 = 11'h6d7 == cnt[10:0] ? $signed(-32'sh70a3) : $signed(_GEN_3799); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3801 = 11'h6d8 == cnt[10:0] ? $signed(-32'sh7049) : $signed(_GEN_3800); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3802 = 11'h6d9 == cnt[10:0] ? $signed(-32'sh6fef) : $signed(_GEN_3801); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3803 = 11'h6da == cnt[10:0] ? $signed(-32'sh6f94) : $signed(_GEN_3802); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3804 = 11'h6db == cnt[10:0] ? $signed(-32'sh6f3a) : $signed(_GEN_3803); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3805 = 11'h6dc == cnt[10:0] ? $signed(-32'sh6edf) : $signed(_GEN_3804); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3806 = 11'h6dd == cnt[10:0] ? $signed(-32'sh6e85) : $signed(_GEN_3805); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3807 = 11'h6de == cnt[10:0] ? $signed(-32'sh6e2a) : $signed(_GEN_3806); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3808 = 11'h6df == cnt[10:0] ? $signed(-32'sh6dcf) : $signed(_GEN_3807); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3809 = 11'h6e0 == cnt[10:0] ? $signed(-32'sh6d74) : $signed(_GEN_3808); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3810 = 11'h6e1 == cnt[10:0] ? $signed(-32'sh6d19) : $signed(_GEN_3809); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3811 = 11'h6e2 == cnt[10:0] ? $signed(-32'sh6cbe) : $signed(_GEN_3810); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3812 = 11'h6e3 == cnt[10:0] ? $signed(-32'sh6c63) : $signed(_GEN_3811); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3813 = 11'h6e4 == cnt[10:0] ? $signed(-32'sh6c08) : $signed(_GEN_3812); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3814 = 11'h6e5 == cnt[10:0] ? $signed(-32'sh6bad) : $signed(_GEN_3813); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3815 = 11'h6e6 == cnt[10:0] ? $signed(-32'sh6b52) : $signed(_GEN_3814); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3816 = 11'h6e7 == cnt[10:0] ? $signed(-32'sh6af6) : $signed(_GEN_3815); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3817 = 11'h6e8 == cnt[10:0] ? $signed(-32'sh6a9b) : $signed(_GEN_3816); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3818 = 11'h6e9 == cnt[10:0] ? $signed(-32'sh6a40) : $signed(_GEN_3817); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3819 = 11'h6ea == cnt[10:0] ? $signed(-32'sh69e4) : $signed(_GEN_3818); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3820 = 11'h6eb == cnt[10:0] ? $signed(-32'sh6989) : $signed(_GEN_3819); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3821 = 11'h6ec == cnt[10:0] ? $signed(-32'sh692d) : $signed(_GEN_3820); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3822 = 11'h6ed == cnt[10:0] ? $signed(-32'sh68d1) : $signed(_GEN_3821); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3823 = 11'h6ee == cnt[10:0] ? $signed(-32'sh6876) : $signed(_GEN_3822); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3824 = 11'h6ef == cnt[10:0] ? $signed(-32'sh681a) : $signed(_GEN_3823); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3825 = 11'h6f0 == cnt[10:0] ? $signed(-32'sh67be) : $signed(_GEN_3824); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3826 = 11'h6f1 == cnt[10:0] ? $signed(-32'sh6762) : $signed(_GEN_3825); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3827 = 11'h6f2 == cnt[10:0] ? $signed(-32'sh6706) : $signed(_GEN_3826); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3828 = 11'h6f3 == cnt[10:0] ? $signed(-32'sh66aa) : $signed(_GEN_3827); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3829 = 11'h6f4 == cnt[10:0] ? $signed(-32'sh664e) : $signed(_GEN_3828); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3830 = 11'h6f5 == cnt[10:0] ? $signed(-32'sh65f2) : $signed(_GEN_3829); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3831 = 11'h6f6 == cnt[10:0] ? $signed(-32'sh6595) : $signed(_GEN_3830); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3832 = 11'h6f7 == cnt[10:0] ? $signed(-32'sh6539) : $signed(_GEN_3831); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3833 = 11'h6f8 == cnt[10:0] ? $signed(-32'sh64dd) : $signed(_GEN_3832); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3834 = 11'h6f9 == cnt[10:0] ? $signed(-32'sh6480) : $signed(_GEN_3833); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3835 = 11'h6fa == cnt[10:0] ? $signed(-32'sh6424) : $signed(_GEN_3834); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3836 = 11'h6fb == cnt[10:0] ? $signed(-32'sh63c7) : $signed(_GEN_3835); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3837 = 11'h6fc == cnt[10:0] ? $signed(-32'sh636b) : $signed(_GEN_3836); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3838 = 11'h6fd == cnt[10:0] ? $signed(-32'sh630e) : $signed(_GEN_3837); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3839 = 11'h6fe == cnt[10:0] ? $signed(-32'sh62b1) : $signed(_GEN_3838); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3840 = 11'h6ff == cnt[10:0] ? $signed(-32'sh6254) : $signed(_GEN_3839); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3841 = 11'h700 == cnt[10:0] ? $signed(-32'sh61f8) : $signed(_GEN_3840); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3842 = 11'h701 == cnt[10:0] ? $signed(-32'sh619b) : $signed(_GEN_3841); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3843 = 11'h702 == cnt[10:0] ? $signed(-32'sh613e) : $signed(_GEN_3842); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3844 = 11'h703 == cnt[10:0] ? $signed(-32'sh60e1) : $signed(_GEN_3843); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3845 = 11'h704 == cnt[10:0] ? $signed(-32'sh6084) : $signed(_GEN_3844); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3846 = 11'h705 == cnt[10:0] ? $signed(-32'sh6026) : $signed(_GEN_3845); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3847 = 11'h706 == cnt[10:0] ? $signed(-32'sh5fc9) : $signed(_GEN_3846); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3848 = 11'h707 == cnt[10:0] ? $signed(-32'sh5f6c) : $signed(_GEN_3847); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3849 = 11'h708 == cnt[10:0] ? $signed(-32'sh5f0f) : $signed(_GEN_3848); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3850 = 11'h709 == cnt[10:0] ? $signed(-32'sh5eb1) : $signed(_GEN_3849); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3851 = 11'h70a == cnt[10:0] ? $signed(-32'sh5e54) : $signed(_GEN_3850); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3852 = 11'h70b == cnt[10:0] ? $signed(-32'sh5df6) : $signed(_GEN_3851); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3853 = 11'h70c == cnt[10:0] ? $signed(-32'sh5d99) : $signed(_GEN_3852); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3854 = 11'h70d == cnt[10:0] ? $signed(-32'sh5d3b) : $signed(_GEN_3853); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3855 = 11'h70e == cnt[10:0] ? $signed(-32'sh5cde) : $signed(_GEN_3854); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3856 = 11'h70f == cnt[10:0] ? $signed(-32'sh5c80) : $signed(_GEN_3855); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3857 = 11'h710 == cnt[10:0] ? $signed(-32'sh5c22) : $signed(_GEN_3856); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3858 = 11'h711 == cnt[10:0] ? $signed(-32'sh5bc4) : $signed(_GEN_3857); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3859 = 11'h712 == cnt[10:0] ? $signed(-32'sh5b66) : $signed(_GEN_3858); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3860 = 11'h713 == cnt[10:0] ? $signed(-32'sh5b08) : $signed(_GEN_3859); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3861 = 11'h714 == cnt[10:0] ? $signed(-32'sh5aaa) : $signed(_GEN_3860); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3862 = 11'h715 == cnt[10:0] ? $signed(-32'sh5a4c) : $signed(_GEN_3861); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3863 = 11'h716 == cnt[10:0] ? $signed(-32'sh59ee) : $signed(_GEN_3862); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3864 = 11'h717 == cnt[10:0] ? $signed(-32'sh5990) : $signed(_GEN_3863); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3865 = 11'h718 == cnt[10:0] ? $signed(-32'sh5932) : $signed(_GEN_3864); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3866 = 11'h719 == cnt[10:0] ? $signed(-32'sh58d4) : $signed(_GEN_3865); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3867 = 11'h71a == cnt[10:0] ? $signed(-32'sh5875) : $signed(_GEN_3866); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3868 = 11'h71b == cnt[10:0] ? $signed(-32'sh5817) : $signed(_GEN_3867); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3869 = 11'h71c == cnt[10:0] ? $signed(-32'sh57b9) : $signed(_GEN_3868); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3870 = 11'h71d == cnt[10:0] ? $signed(-32'sh575a) : $signed(_GEN_3869); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3871 = 11'h71e == cnt[10:0] ? $signed(-32'sh56fc) : $signed(_GEN_3870); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3872 = 11'h71f == cnt[10:0] ? $signed(-32'sh569d) : $signed(_GEN_3871); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3873 = 11'h720 == cnt[10:0] ? $signed(-32'sh563e) : $signed(_GEN_3872); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3874 = 11'h721 == cnt[10:0] ? $signed(-32'sh55e0) : $signed(_GEN_3873); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3875 = 11'h722 == cnt[10:0] ? $signed(-32'sh5581) : $signed(_GEN_3874); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3876 = 11'h723 == cnt[10:0] ? $signed(-32'sh5522) : $signed(_GEN_3875); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3877 = 11'h724 == cnt[10:0] ? $signed(-32'sh54c3) : $signed(_GEN_3876); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3878 = 11'h725 == cnt[10:0] ? $signed(-32'sh5464) : $signed(_GEN_3877); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3879 = 11'h726 == cnt[10:0] ? $signed(-32'sh5406) : $signed(_GEN_3878); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3880 = 11'h727 == cnt[10:0] ? $signed(-32'sh53a7) : $signed(_GEN_3879); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3881 = 11'h728 == cnt[10:0] ? $signed(-32'sh5348) : $signed(_GEN_3880); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3882 = 11'h729 == cnt[10:0] ? $signed(-32'sh52e8) : $signed(_GEN_3881); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3883 = 11'h72a == cnt[10:0] ? $signed(-32'sh5289) : $signed(_GEN_3882); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3884 = 11'h72b == cnt[10:0] ? $signed(-32'sh522a) : $signed(_GEN_3883); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3885 = 11'h72c == cnt[10:0] ? $signed(-32'sh51cb) : $signed(_GEN_3884); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3886 = 11'h72d == cnt[10:0] ? $signed(-32'sh516c) : $signed(_GEN_3885); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3887 = 11'h72e == cnt[10:0] ? $signed(-32'sh510c) : $signed(_GEN_3886); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3888 = 11'h72f == cnt[10:0] ? $signed(-32'sh50ad) : $signed(_GEN_3887); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3889 = 11'h730 == cnt[10:0] ? $signed(-32'sh504d) : $signed(_GEN_3888); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3890 = 11'h731 == cnt[10:0] ? $signed(-32'sh4fee) : $signed(_GEN_3889); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3891 = 11'h732 == cnt[10:0] ? $signed(-32'sh4f8e) : $signed(_GEN_3890); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3892 = 11'h733 == cnt[10:0] ? $signed(-32'sh4f2f) : $signed(_GEN_3891); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3893 = 11'h734 == cnt[10:0] ? $signed(-32'sh4ecf) : $signed(_GEN_3892); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3894 = 11'h735 == cnt[10:0] ? $signed(-32'sh4e70) : $signed(_GEN_3893); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3895 = 11'h736 == cnt[10:0] ? $signed(-32'sh4e10) : $signed(_GEN_3894); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3896 = 11'h737 == cnt[10:0] ? $signed(-32'sh4db0) : $signed(_GEN_3895); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3897 = 11'h738 == cnt[10:0] ? $signed(-32'sh4d50) : $signed(_GEN_3896); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3898 = 11'h739 == cnt[10:0] ? $signed(-32'sh4cf0) : $signed(_GEN_3897); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3899 = 11'h73a == cnt[10:0] ? $signed(-32'sh4c90) : $signed(_GEN_3898); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3900 = 11'h73b == cnt[10:0] ? $signed(-32'sh4c31) : $signed(_GEN_3899); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3901 = 11'h73c == cnt[10:0] ? $signed(-32'sh4bd1) : $signed(_GEN_3900); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3902 = 11'h73d == cnt[10:0] ? $signed(-32'sh4b71) : $signed(_GEN_3901); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3903 = 11'h73e == cnt[10:0] ? $signed(-32'sh4b10) : $signed(_GEN_3902); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3904 = 11'h73f == cnt[10:0] ? $signed(-32'sh4ab0) : $signed(_GEN_3903); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3905 = 11'h740 == cnt[10:0] ? $signed(-32'sh4a50) : $signed(_GEN_3904); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3906 = 11'h741 == cnt[10:0] ? $signed(-32'sh49f0) : $signed(_GEN_3905); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3907 = 11'h742 == cnt[10:0] ? $signed(-32'sh4990) : $signed(_GEN_3906); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3908 = 11'h743 == cnt[10:0] ? $signed(-32'sh492f) : $signed(_GEN_3907); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3909 = 11'h744 == cnt[10:0] ? $signed(-32'sh48cf) : $signed(_GEN_3908); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3910 = 11'h745 == cnt[10:0] ? $signed(-32'sh486f) : $signed(_GEN_3909); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3911 = 11'h746 == cnt[10:0] ? $signed(-32'sh480e) : $signed(_GEN_3910); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3912 = 11'h747 == cnt[10:0] ? $signed(-32'sh47ae) : $signed(_GEN_3911); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3913 = 11'h748 == cnt[10:0] ? $signed(-32'sh474d) : $signed(_GEN_3912); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3914 = 11'h749 == cnt[10:0] ? $signed(-32'sh46ec) : $signed(_GEN_3913); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3915 = 11'h74a == cnt[10:0] ? $signed(-32'sh468c) : $signed(_GEN_3914); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3916 = 11'h74b == cnt[10:0] ? $signed(-32'sh462b) : $signed(_GEN_3915); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3917 = 11'h74c == cnt[10:0] ? $signed(-32'sh45cb) : $signed(_GEN_3916); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3918 = 11'h74d == cnt[10:0] ? $signed(-32'sh456a) : $signed(_GEN_3917); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3919 = 11'h74e == cnt[10:0] ? $signed(-32'sh4509) : $signed(_GEN_3918); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3920 = 11'h74f == cnt[10:0] ? $signed(-32'sh44a8) : $signed(_GEN_3919); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3921 = 11'h750 == cnt[10:0] ? $signed(-32'sh4447) : $signed(_GEN_3920); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3922 = 11'h751 == cnt[10:0] ? $signed(-32'sh43e6) : $signed(_GEN_3921); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3923 = 11'h752 == cnt[10:0] ? $signed(-32'sh4385) : $signed(_GEN_3922); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3924 = 11'h753 == cnt[10:0] ? $signed(-32'sh4324) : $signed(_GEN_3923); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3925 = 11'h754 == cnt[10:0] ? $signed(-32'sh42c3) : $signed(_GEN_3924); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3926 = 11'h755 == cnt[10:0] ? $signed(-32'sh4262) : $signed(_GEN_3925); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3927 = 11'h756 == cnt[10:0] ? $signed(-32'sh4201) : $signed(_GEN_3926); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3928 = 11'h757 == cnt[10:0] ? $signed(-32'sh41a0) : $signed(_GEN_3927); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3929 = 11'h758 == cnt[10:0] ? $signed(-32'sh413f) : $signed(_GEN_3928); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3930 = 11'h759 == cnt[10:0] ? $signed(-32'sh40de) : $signed(_GEN_3929); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3931 = 11'h75a == cnt[10:0] ? $signed(-32'sh407c) : $signed(_GEN_3930); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3932 = 11'h75b == cnt[10:0] ? $signed(-32'sh401b) : $signed(_GEN_3931); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3933 = 11'h75c == cnt[10:0] ? $signed(-32'sh3fba) : $signed(_GEN_3932); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3934 = 11'h75d == cnt[10:0] ? $signed(-32'sh3f58) : $signed(_GEN_3933); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3935 = 11'h75e == cnt[10:0] ? $signed(-32'sh3ef7) : $signed(_GEN_3934); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3936 = 11'h75f == cnt[10:0] ? $signed(-32'sh3e95) : $signed(_GEN_3935); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3937 = 11'h760 == cnt[10:0] ? $signed(-32'sh3e34) : $signed(_GEN_3936); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3938 = 11'h761 == cnt[10:0] ? $signed(-32'sh3dd2) : $signed(_GEN_3937); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3939 = 11'h762 == cnt[10:0] ? $signed(-32'sh3d71) : $signed(_GEN_3938); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3940 = 11'h763 == cnt[10:0] ? $signed(-32'sh3d0f) : $signed(_GEN_3939); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3941 = 11'h764 == cnt[10:0] ? $signed(-32'sh3cae) : $signed(_GEN_3940); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3942 = 11'h765 == cnt[10:0] ? $signed(-32'sh3c4c) : $signed(_GEN_3941); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3943 = 11'h766 == cnt[10:0] ? $signed(-32'sh3bea) : $signed(_GEN_3942); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3944 = 11'h767 == cnt[10:0] ? $signed(-32'sh3b88) : $signed(_GEN_3943); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3945 = 11'h768 == cnt[10:0] ? $signed(-32'sh3b27) : $signed(_GEN_3944); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3946 = 11'h769 == cnt[10:0] ? $signed(-32'sh3ac5) : $signed(_GEN_3945); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3947 = 11'h76a == cnt[10:0] ? $signed(-32'sh3a63) : $signed(_GEN_3946); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3948 = 11'h76b == cnt[10:0] ? $signed(-32'sh3a01) : $signed(_GEN_3947); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3949 = 11'h76c == cnt[10:0] ? $signed(-32'sh399f) : $signed(_GEN_3948); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3950 = 11'h76d == cnt[10:0] ? $signed(-32'sh393d) : $signed(_GEN_3949); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3951 = 11'h76e == cnt[10:0] ? $signed(-32'sh38db) : $signed(_GEN_3950); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3952 = 11'h76f == cnt[10:0] ? $signed(-32'sh3879) : $signed(_GEN_3951); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3953 = 11'h770 == cnt[10:0] ? $signed(-32'sh3817) : $signed(_GEN_3952); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3954 = 11'h771 == cnt[10:0] ? $signed(-32'sh37b5) : $signed(_GEN_3953); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3955 = 11'h772 == cnt[10:0] ? $signed(-32'sh3753) : $signed(_GEN_3954); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3956 = 11'h773 == cnt[10:0] ? $signed(-32'sh36f1) : $signed(_GEN_3955); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3957 = 11'h774 == cnt[10:0] ? $signed(-32'sh368e) : $signed(_GEN_3956); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3958 = 11'h775 == cnt[10:0] ? $signed(-32'sh362c) : $signed(_GEN_3957); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3959 = 11'h776 == cnt[10:0] ? $signed(-32'sh35ca) : $signed(_GEN_3958); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3960 = 11'h777 == cnt[10:0] ? $signed(-32'sh3568) : $signed(_GEN_3959); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3961 = 11'h778 == cnt[10:0] ? $signed(-32'sh3505) : $signed(_GEN_3960); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3962 = 11'h779 == cnt[10:0] ? $signed(-32'sh34a3) : $signed(_GEN_3961); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3963 = 11'h77a == cnt[10:0] ? $signed(-32'sh3440) : $signed(_GEN_3962); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3964 = 11'h77b == cnt[10:0] ? $signed(-32'sh33de) : $signed(_GEN_3963); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3965 = 11'h77c == cnt[10:0] ? $signed(-32'sh337c) : $signed(_GEN_3964); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3966 = 11'h77d == cnt[10:0] ? $signed(-32'sh3319) : $signed(_GEN_3965); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3967 = 11'h77e == cnt[10:0] ? $signed(-32'sh32b7) : $signed(_GEN_3966); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3968 = 11'h77f == cnt[10:0] ? $signed(-32'sh3254) : $signed(_GEN_3967); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3969 = 11'h780 == cnt[10:0] ? $signed(-32'sh31f1) : $signed(_GEN_3968); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3970 = 11'h781 == cnt[10:0] ? $signed(-32'sh318f) : $signed(_GEN_3969); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3971 = 11'h782 == cnt[10:0] ? $signed(-32'sh312c) : $signed(_GEN_3970); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3972 = 11'h783 == cnt[10:0] ? $signed(-32'sh30ca) : $signed(_GEN_3971); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3973 = 11'h784 == cnt[10:0] ? $signed(-32'sh3067) : $signed(_GEN_3972); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3974 = 11'h785 == cnt[10:0] ? $signed(-32'sh3004) : $signed(_GEN_3973); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3975 = 11'h786 == cnt[10:0] ? $signed(-32'sh2fa1) : $signed(_GEN_3974); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3976 = 11'h787 == cnt[10:0] ? $signed(-32'sh2f3f) : $signed(_GEN_3975); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3977 = 11'h788 == cnt[10:0] ? $signed(-32'sh2edc) : $signed(_GEN_3976); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3978 = 11'h789 == cnt[10:0] ? $signed(-32'sh2e79) : $signed(_GEN_3977); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3979 = 11'h78a == cnt[10:0] ? $signed(-32'sh2e16) : $signed(_GEN_3978); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3980 = 11'h78b == cnt[10:0] ? $signed(-32'sh2db3) : $signed(_GEN_3979); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3981 = 11'h78c == cnt[10:0] ? $signed(-32'sh2d50) : $signed(_GEN_3980); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3982 = 11'h78d == cnt[10:0] ? $signed(-32'sh2ced) : $signed(_GEN_3981); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3983 = 11'h78e == cnt[10:0] ? $signed(-32'sh2c8a) : $signed(_GEN_3982); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3984 = 11'h78f == cnt[10:0] ? $signed(-32'sh2c27) : $signed(_GEN_3983); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3985 = 11'h790 == cnt[10:0] ? $signed(-32'sh2bc4) : $signed(_GEN_3984); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3986 = 11'h791 == cnt[10:0] ? $signed(-32'sh2b61) : $signed(_GEN_3985); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3987 = 11'h792 == cnt[10:0] ? $signed(-32'sh2afe) : $signed(_GEN_3986); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3988 = 11'h793 == cnt[10:0] ? $signed(-32'sh2a9b) : $signed(_GEN_3987); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3989 = 11'h794 == cnt[10:0] ? $signed(-32'sh2a38) : $signed(_GEN_3988); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3990 = 11'h795 == cnt[10:0] ? $signed(-32'sh29d5) : $signed(_GEN_3989); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3991 = 11'h796 == cnt[10:0] ? $signed(-32'sh2971) : $signed(_GEN_3990); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3992 = 11'h797 == cnt[10:0] ? $signed(-32'sh290e) : $signed(_GEN_3991); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3993 = 11'h798 == cnt[10:0] ? $signed(-32'sh28ab) : $signed(_GEN_3992); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3994 = 11'h799 == cnt[10:0] ? $signed(-32'sh2848) : $signed(_GEN_3993); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3995 = 11'h79a == cnt[10:0] ? $signed(-32'sh27e4) : $signed(_GEN_3994); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3996 = 11'h79b == cnt[10:0] ? $signed(-32'sh2781) : $signed(_GEN_3995); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3997 = 11'h79c == cnt[10:0] ? $signed(-32'sh271e) : $signed(_GEN_3996); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3998 = 11'h79d == cnt[10:0] ? $signed(-32'sh26ba) : $signed(_GEN_3997); // @[FFT.scala 35:12]
  wire [31:0] _GEN_3999 = 11'h79e == cnt[10:0] ? $signed(-32'sh2657) : $signed(_GEN_3998); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4000 = 11'h79f == cnt[10:0] ? $signed(-32'sh25f4) : $signed(_GEN_3999); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4001 = 11'h7a0 == cnt[10:0] ? $signed(-32'sh2590) : $signed(_GEN_4000); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4002 = 11'h7a1 == cnt[10:0] ? $signed(-32'sh252d) : $signed(_GEN_4001); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4003 = 11'h7a2 == cnt[10:0] ? $signed(-32'sh24c9) : $signed(_GEN_4002); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4004 = 11'h7a3 == cnt[10:0] ? $signed(-32'sh2466) : $signed(_GEN_4003); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4005 = 11'h7a4 == cnt[10:0] ? $signed(-32'sh2402) : $signed(_GEN_4004); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4006 = 11'h7a5 == cnt[10:0] ? $signed(-32'sh239f) : $signed(_GEN_4005); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4007 = 11'h7a6 == cnt[10:0] ? $signed(-32'sh233b) : $signed(_GEN_4006); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4008 = 11'h7a7 == cnt[10:0] ? $signed(-32'sh22d7) : $signed(_GEN_4007); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4009 = 11'h7a8 == cnt[10:0] ? $signed(-32'sh2274) : $signed(_GEN_4008); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4010 = 11'h7a9 == cnt[10:0] ? $signed(-32'sh2210) : $signed(_GEN_4009); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4011 = 11'h7aa == cnt[10:0] ? $signed(-32'sh21ad) : $signed(_GEN_4010); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4012 = 11'h7ab == cnt[10:0] ? $signed(-32'sh2149) : $signed(_GEN_4011); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4013 = 11'h7ac == cnt[10:0] ? $signed(-32'sh20e5) : $signed(_GEN_4012); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4014 = 11'h7ad == cnt[10:0] ? $signed(-32'sh2082) : $signed(_GEN_4013); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4015 = 11'h7ae == cnt[10:0] ? $signed(-32'sh201e) : $signed(_GEN_4014); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4016 = 11'h7af == cnt[10:0] ? $signed(-32'sh1fba) : $signed(_GEN_4015); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4017 = 11'h7b0 == cnt[10:0] ? $signed(-32'sh1f56) : $signed(_GEN_4016); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4018 = 11'h7b1 == cnt[10:0] ? $signed(-32'sh1ef3) : $signed(_GEN_4017); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4019 = 11'h7b2 == cnt[10:0] ? $signed(-32'sh1e8f) : $signed(_GEN_4018); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4020 = 11'h7b3 == cnt[10:0] ? $signed(-32'sh1e2b) : $signed(_GEN_4019); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4021 = 11'h7b4 == cnt[10:0] ? $signed(-32'sh1dc7) : $signed(_GEN_4020); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4022 = 11'h7b5 == cnt[10:0] ? $signed(-32'sh1d63) : $signed(_GEN_4021); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4023 = 11'h7b6 == cnt[10:0] ? $signed(-32'sh1cff) : $signed(_GEN_4022); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4024 = 11'h7b7 == cnt[10:0] ? $signed(-32'sh1c9b) : $signed(_GEN_4023); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4025 = 11'h7b8 == cnt[10:0] ? $signed(-32'sh1c38) : $signed(_GEN_4024); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4026 = 11'h7b9 == cnt[10:0] ? $signed(-32'sh1bd4) : $signed(_GEN_4025); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4027 = 11'h7ba == cnt[10:0] ? $signed(-32'sh1b70) : $signed(_GEN_4026); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4028 = 11'h7bb == cnt[10:0] ? $signed(-32'sh1b0c) : $signed(_GEN_4027); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4029 = 11'h7bc == cnt[10:0] ? $signed(-32'sh1aa8) : $signed(_GEN_4028); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4030 = 11'h7bd == cnt[10:0] ? $signed(-32'sh1a44) : $signed(_GEN_4029); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4031 = 11'h7be == cnt[10:0] ? $signed(-32'sh19e0) : $signed(_GEN_4030); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4032 = 11'h7bf == cnt[10:0] ? $signed(-32'sh197c) : $signed(_GEN_4031); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4033 = 11'h7c0 == cnt[10:0] ? $signed(-32'sh1918) : $signed(_GEN_4032); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4034 = 11'h7c1 == cnt[10:0] ? $signed(-32'sh18b4) : $signed(_GEN_4033); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4035 = 11'h7c2 == cnt[10:0] ? $signed(-32'sh1850) : $signed(_GEN_4034); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4036 = 11'h7c3 == cnt[10:0] ? $signed(-32'sh17eb) : $signed(_GEN_4035); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4037 = 11'h7c4 == cnt[10:0] ? $signed(-32'sh1787) : $signed(_GEN_4036); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4038 = 11'h7c5 == cnt[10:0] ? $signed(-32'sh1723) : $signed(_GEN_4037); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4039 = 11'h7c6 == cnt[10:0] ? $signed(-32'sh16bf) : $signed(_GEN_4038); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4040 = 11'h7c7 == cnt[10:0] ? $signed(-32'sh165b) : $signed(_GEN_4039); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4041 = 11'h7c8 == cnt[10:0] ? $signed(-32'sh15f7) : $signed(_GEN_4040); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4042 = 11'h7c9 == cnt[10:0] ? $signed(-32'sh1593) : $signed(_GEN_4041); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4043 = 11'h7ca == cnt[10:0] ? $signed(-32'sh152e) : $signed(_GEN_4042); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4044 = 11'h7cb == cnt[10:0] ? $signed(-32'sh14ca) : $signed(_GEN_4043); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4045 = 11'h7cc == cnt[10:0] ? $signed(-32'sh1466) : $signed(_GEN_4044); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4046 = 11'h7cd == cnt[10:0] ? $signed(-32'sh1402) : $signed(_GEN_4045); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4047 = 11'h7ce == cnt[10:0] ? $signed(-32'sh139e) : $signed(_GEN_4046); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4048 = 11'h7cf == cnt[10:0] ? $signed(-32'sh1339) : $signed(_GEN_4047); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4049 = 11'h7d0 == cnt[10:0] ? $signed(-32'sh12d5) : $signed(_GEN_4048); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4050 = 11'h7d1 == cnt[10:0] ? $signed(-32'sh1271) : $signed(_GEN_4049); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4051 = 11'h7d2 == cnt[10:0] ? $signed(-32'sh120d) : $signed(_GEN_4050); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4052 = 11'h7d3 == cnt[10:0] ? $signed(-32'sh11a8) : $signed(_GEN_4051); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4053 = 11'h7d4 == cnt[10:0] ? $signed(-32'sh1144) : $signed(_GEN_4052); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4054 = 11'h7d5 == cnt[10:0] ? $signed(-32'sh10e0) : $signed(_GEN_4053); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4055 = 11'h7d6 == cnt[10:0] ? $signed(-32'sh107b) : $signed(_GEN_4054); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4056 = 11'h7d7 == cnt[10:0] ? $signed(-32'sh1017) : $signed(_GEN_4055); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4057 = 11'h7d8 == cnt[10:0] ? $signed(-32'shfb3) : $signed(_GEN_4056); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4058 = 11'h7d9 == cnt[10:0] ? $signed(-32'shf4e) : $signed(_GEN_4057); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4059 = 11'h7da == cnt[10:0] ? $signed(-32'sheea) : $signed(_GEN_4058); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4060 = 11'h7db == cnt[10:0] ? $signed(-32'she86) : $signed(_GEN_4059); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4061 = 11'h7dc == cnt[10:0] ? $signed(-32'she21) : $signed(_GEN_4060); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4062 = 11'h7dd == cnt[10:0] ? $signed(-32'shdbd) : $signed(_GEN_4061); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4063 = 11'h7de == cnt[10:0] ? $signed(-32'shd59) : $signed(_GEN_4062); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4064 = 11'h7df == cnt[10:0] ? $signed(-32'shcf4) : $signed(_GEN_4063); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4065 = 11'h7e0 == cnt[10:0] ? $signed(-32'shc90) : $signed(_GEN_4064); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4066 = 11'h7e1 == cnt[10:0] ? $signed(-32'shc2b) : $signed(_GEN_4065); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4067 = 11'h7e2 == cnt[10:0] ? $signed(-32'shbc7) : $signed(_GEN_4066); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4068 = 11'h7e3 == cnt[10:0] ? $signed(-32'shb62) : $signed(_GEN_4067); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4069 = 11'h7e4 == cnt[10:0] ? $signed(-32'shafe) : $signed(_GEN_4068); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4070 = 11'h7e5 == cnt[10:0] ? $signed(-32'sha9a) : $signed(_GEN_4069); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4071 = 11'h7e6 == cnt[10:0] ? $signed(-32'sha35) : $signed(_GEN_4070); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4072 = 11'h7e7 == cnt[10:0] ? $signed(-32'sh9d1) : $signed(_GEN_4071); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4073 = 11'h7e8 == cnt[10:0] ? $signed(-32'sh96c) : $signed(_GEN_4072); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4074 = 11'h7e9 == cnt[10:0] ? $signed(-32'sh908) : $signed(_GEN_4073); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4075 = 11'h7ea == cnt[10:0] ? $signed(-32'sh8a3) : $signed(_GEN_4074); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4076 = 11'h7eb == cnt[10:0] ? $signed(-32'sh83f) : $signed(_GEN_4075); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4077 = 11'h7ec == cnt[10:0] ? $signed(-32'sh7da) : $signed(_GEN_4076); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4078 = 11'h7ed == cnt[10:0] ? $signed(-32'sh776) : $signed(_GEN_4077); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4079 = 11'h7ee == cnt[10:0] ? $signed(-32'sh711) : $signed(_GEN_4078); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4080 = 11'h7ef == cnt[10:0] ? $signed(-32'sh6ad) : $signed(_GEN_4079); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4081 = 11'h7f0 == cnt[10:0] ? $signed(-32'sh648) : $signed(_GEN_4080); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4082 = 11'h7f1 == cnt[10:0] ? $signed(-32'sh5e4) : $signed(_GEN_4081); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4083 = 11'h7f2 == cnt[10:0] ? $signed(-32'sh57f) : $signed(_GEN_4082); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4084 = 11'h7f3 == cnt[10:0] ? $signed(-32'sh51b) : $signed(_GEN_4083); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4085 = 11'h7f4 == cnt[10:0] ? $signed(-32'sh4b6) : $signed(_GEN_4084); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4086 = 11'h7f5 == cnt[10:0] ? $signed(-32'sh452) : $signed(_GEN_4085); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4087 = 11'h7f6 == cnt[10:0] ? $signed(-32'sh3ed) : $signed(_GEN_4086); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4088 = 11'h7f7 == cnt[10:0] ? $signed(-32'sh389) : $signed(_GEN_4087); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4089 = 11'h7f8 == cnt[10:0] ? $signed(-32'sh324) : $signed(_GEN_4088); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4090 = 11'h7f9 == cnt[10:0] ? $signed(-32'sh2c0) : $signed(_GEN_4089); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4091 = 11'h7fa == cnt[10:0] ? $signed(-32'sh25b) : $signed(_GEN_4090); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4092 = 11'h7fb == cnt[10:0] ? $signed(-32'sh1f7) : $signed(_GEN_4091); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4093 = 11'h7fc == cnt[10:0] ? $signed(-32'sh192) : $signed(_GEN_4092); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4094 = 11'h7fd == cnt[10:0] ? $signed(-32'sh12e) : $signed(_GEN_4093); // @[FFT.scala 35:12]
  wire [31:0] _GEN_4095 = 11'h7fe == cnt[10:0] ? $signed(-32'shc9) : $signed(_GEN_4094); // @[FFT.scala 35:12]
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_763;
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_764;
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_765;
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_766;
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_767;
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_768;
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg [31:0] _T_674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg [31:0] _T_674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1025;
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1026;
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1027;
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1028;
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1029;
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1030;
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1031;
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1032;
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1033;
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1034;
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1035;
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1036;
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1037;
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1038;
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1039;
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1040;
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1041;
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1042;
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1043;
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1044;
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1045;
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1046;
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1047;
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1048;
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1049;
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1050;
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1051;
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1052;
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1053;
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1054;
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1055;
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1056;
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1057;
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1058;
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1059;
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1060;
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1061;
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1062;
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1063;
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1064;
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1065;
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1066;
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1067;
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1068;
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1069;
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1070;
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1071;
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1072;
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1073;
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1074;
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1075;
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1076;
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1077;
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1078;
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1079;
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1080;
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1081;
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1082;
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1083;
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1084;
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1085;
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1086;
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1087;
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1088;
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1089;
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1090;
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1091;
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1092;
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1093;
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1094;
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1095;
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1096;
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1097;
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1098;
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1099;
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1100;
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1101;
  reg [31:0] _T_739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1102;
  reg [31:0] _T_739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1103;
  reg [31:0] _T_740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1104;
  reg [31:0] _T_740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1105;
  reg [31:0] _T_741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1106;
  reg [31:0] _T_741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1107;
  reg [31:0] _T_742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1108;
  reg [31:0] _T_742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1109;
  reg [31:0] _T_743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1110;
  reg [31:0] _T_743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1111;
  reg [31:0] _T_744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1112;
  reg [31:0] _T_744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1113;
  reg [31:0] _T_745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1114;
  reg [31:0] _T_745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1115;
  reg [31:0] _T_746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1116;
  reg [31:0] _T_746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1117;
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1118;
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1119;
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1120;
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1121;
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1122;
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1123;
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1124;
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1125;
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1126;
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1127;
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1128;
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1129;
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1130;
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1131;
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1132;
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1133;
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1134;
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1135;
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1136;
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1137;
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1138;
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1139;
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1140;
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1141;
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1142;
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1143;
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1144;
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1145;
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1146;
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1147;
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1148;
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1149;
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1150;
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1151;
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1152;
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1153;
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1154;
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1155;
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1156;
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1157;
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1158;
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1159;
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1160;
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1161;
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1162;
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1163;
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1164;
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1165;
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1166;
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1167;
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1168;
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1169;
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1170;
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1171;
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1172;
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1173;
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1174;
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1175;
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1176;
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1177;
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1178;
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1179;
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1180;
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1181;
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1182;
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1183;
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1184;
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1185;
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1186;
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1187;
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1188;
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1189;
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1190;
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1191;
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1192;
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1193;
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1194;
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1195;
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1196;
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1197;
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1198;
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1199;
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1200;
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1201;
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1202;
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1203;
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1204;
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1205;
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1206;
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1207;
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1208;
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1209;
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1210;
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1211;
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1212;
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1213;
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1214;
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1215;
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1216;
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1217;
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1218;
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1219;
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1220;
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1221;
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1222;
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1223;
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1224;
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1225;
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1226;
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1227;
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1228;
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1229;
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1230;
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1231;
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1232;
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1233;
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1234;
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1235;
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1236;
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1237;
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1238;
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1239;
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1240;
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1241;
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1242;
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1243;
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1244;
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1245;
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1246;
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1247;
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1248;
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1249;
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1250;
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1251;
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1252;
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1253;
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1254;
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1255;
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1256;
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1257;
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1258;
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1259;
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1260;
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1261;
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1262;
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1263;
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1264;
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1265;
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1266;
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1267;
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1268;
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1269;
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1270;
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1271;
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1272;
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1273;
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1274;
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1275;
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1276;
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1277;
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1278;
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1279;
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1280;
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1281;
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1282;
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1283;
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1284;
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1285;
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1286;
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1287;
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1288;
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1289;
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1290;
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1291;
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1292;
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1293;
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1294;
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1295;
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1296;
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1297;
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1298;
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1299;
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1300;
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1301;
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1302;
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1303;
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1304;
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1305;
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1306;
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1307;
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1308;
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1309;
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1310;
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1311;
  reg [31:0] _T_844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1312;
  reg [31:0] _T_844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1313;
  reg [31:0] _T_845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1314;
  reg [31:0] _T_845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1315;
  reg [31:0] _T_846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1316;
  reg [31:0] _T_846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1317;
  reg [31:0] _T_847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1318;
  reg [31:0] _T_847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1319;
  reg [31:0] _T_848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1320;
  reg [31:0] _T_848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1321;
  reg [31:0] _T_849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1322;
  reg [31:0] _T_849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1323;
  reg [31:0] _T_850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1324;
  reg [31:0] _T_850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1325;
  reg [31:0] _T_851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1326;
  reg [31:0] _T_851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1327;
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1328;
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1329;
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1330;
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1331;
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1332;
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1333;
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1334;
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1335;
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1336;
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1337;
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1338;
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1339;
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1340;
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1341;
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1342;
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1343;
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1344;
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1345;
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1346;
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1347;
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1348;
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1349;
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1350;
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1351;
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1352;
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1353;
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1354;
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1355;
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1356;
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1357;
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1358;
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1359;
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1360;
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1361;
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1362;
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1363;
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1364;
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1365;
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1366;
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1367;
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1368;
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1369;
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1370;
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1371;
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1372;
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1373;
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1374;
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1375;
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1376;
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1377;
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1378;
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1379;
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1380;
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1381;
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1382;
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1383;
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1384;
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1385;
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1386;
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1387;
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1388;
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1389;
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1390;
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1391;
  reg [31:0] _T_884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1392;
  reg [31:0] _T_884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1393;
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1394;
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1395;
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1396;
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1397;
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1398;
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1399;
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1400;
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1401;
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1402;
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1403;
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1404;
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1405;
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1406;
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1407;
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1408;
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1409;
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1410;
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1411;
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1412;
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1413;
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1414;
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1415;
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1416;
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1417;
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1418;
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1419;
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1420;
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1421;
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1422;
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1423;
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1424;
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1425;
  reg [31:0] _T_901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1426;
  reg [31:0] _T_901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1427;
  reg [31:0] _T_902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1428;
  reg [31:0] _T_902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1429;
  reg [31:0] _T_903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1430;
  reg [31:0] _T_903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1431;
  reg [31:0] _T_904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1432;
  reg [31:0] _T_904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1433;
  reg [31:0] _T_905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1434;
  reg [31:0] _T_905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1435;
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1436;
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1437;
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1438;
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1439;
  reg [31:0] _T_908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1440;
  reg [31:0] _T_908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1441;
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1442;
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1443;
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1444;
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1445;
  reg [31:0] _T_911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1446;
  reg [31:0] _T_911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1447;
  reg [31:0] _T_912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1448;
  reg [31:0] _T_912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1449;
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1450;
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1451;
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1452;
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1453;
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1454;
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1455;
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1456;
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1457;
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1458;
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1459;
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1460;
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1461;
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1462;
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1463;
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1464;
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1465;
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1466;
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1467;
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1468;
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1469;
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1470;
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1471;
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1472;
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1473;
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1474;
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1475;
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1476;
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1477;
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1478;
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1479;
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1480;
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1481;
  reg [31:0] _T_929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1482;
  reg [31:0] _T_929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1483;
  reg [31:0] _T_930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1484;
  reg [31:0] _T_930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1485;
  reg [31:0] _T_931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1486;
  reg [31:0] _T_931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1487;
  reg [31:0] _T_932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1488;
  reg [31:0] _T_932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1489;
  reg [31:0] _T_933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1490;
  reg [31:0] _T_933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1491;
  reg [31:0] _T_934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1492;
  reg [31:0] _T_934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1493;
  reg [31:0] _T_935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1494;
  reg [31:0] _T_935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1495;
  reg [31:0] _T_936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1496;
  reg [31:0] _T_936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1497;
  reg [31:0] _T_937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1498;
  reg [31:0] _T_937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1499;
  reg [31:0] _T_938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1500;
  reg [31:0] _T_938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1501;
  reg [31:0] _T_939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1502;
  reg [31:0] _T_939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1503;
  reg [31:0] _T_940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1504;
  reg [31:0] _T_940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1505;
  reg [31:0] _T_941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1506;
  reg [31:0] _T_941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1507;
  reg [31:0] _T_942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1508;
  reg [31:0] _T_942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1509;
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1510;
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1511;
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1512;
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1513;
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1514;
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1515;
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1516;
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1517;
  reg [31:0] _T_947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1518;
  reg [31:0] _T_947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1519;
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1520;
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1521;
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1522;
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1523;
  reg [31:0] _T_950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1524;
  reg [31:0] _T_950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1525;
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1526;
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1527;
  reg [31:0] _T_952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1528;
  reg [31:0] _T_952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1529;
  reg [31:0] _T_953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1530;
  reg [31:0] _T_953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1531;
  reg [31:0] _T_954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1532;
  reg [31:0] _T_954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1533;
  reg [31:0] _T_955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1534;
  reg [31:0] _T_955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1535;
  reg [31:0] _T_956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1536;
  reg [31:0] _T_956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1537;
  reg [31:0] _T_957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1538;
  reg [31:0] _T_957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1539;
  reg [31:0] _T_958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1540;
  reg [31:0] _T_958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1541;
  reg [31:0] _T_959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1542;
  reg [31:0] _T_959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1543;
  reg [31:0] _T_960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1544;
  reg [31:0] _T_960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1545;
  reg [31:0] _T_961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1546;
  reg [31:0] _T_961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1547;
  reg [31:0] _T_962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1548;
  reg [31:0] _T_962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1549;
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1550;
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1551;
  reg [31:0] _T_964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1552;
  reg [31:0] _T_964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1553;
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1554;
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1555;
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1556;
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1557;
  reg [31:0] _T_967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1558;
  reg [31:0] _T_967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1559;
  reg [31:0] _T_968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1560;
  reg [31:0] _T_968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1561;
  reg [31:0] _T_969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1562;
  reg [31:0] _T_969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1563;
  reg [31:0] _T_970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1564;
  reg [31:0] _T_970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1565;
  reg [31:0] _T_971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1566;
  reg [31:0] _T_971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1567;
  reg [31:0] _T_972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1568;
  reg [31:0] _T_972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1569;
  reg [31:0] _T_973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1570;
  reg [31:0] _T_973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1571;
  reg [31:0] _T_974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1572;
  reg [31:0] _T_974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1573;
  reg [31:0] _T_975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1574;
  reg [31:0] _T_975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1575;
  reg [31:0] _T_976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1576;
  reg [31:0] _T_976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1577;
  reg [31:0] _T_977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1578;
  reg [31:0] _T_977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1579;
  reg [31:0] _T_978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1580;
  reg [31:0] _T_978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1581;
  reg [31:0] _T_979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1582;
  reg [31:0] _T_979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1583;
  reg [31:0] _T_980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1584;
  reg [31:0] _T_980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1585;
  reg [31:0] _T_981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1586;
  reg [31:0] _T_981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1587;
  reg [31:0] _T_982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1588;
  reg [31:0] _T_982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1589;
  reg [31:0] _T_983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1590;
  reg [31:0] _T_983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1591;
  reg [31:0] _T_984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1592;
  reg [31:0] _T_984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1593;
  reg [31:0] _T_985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1594;
  reg [31:0] _T_985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1595;
  reg [31:0] _T_986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1596;
  reg [31:0] _T_986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1597;
  reg [31:0] _T_987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1598;
  reg [31:0] _T_987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1599;
  reg [31:0] _T_988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1600;
  reg [31:0] _T_988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1601;
  reg [31:0] _T_989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1602;
  reg [31:0] _T_989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1603;
  reg [31:0] _T_990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1604;
  reg [31:0] _T_990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1605;
  reg [31:0] _T_991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1606;
  reg [31:0] _T_991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1607;
  reg [31:0] _T_992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1608;
  reg [31:0] _T_992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1609;
  reg [31:0] _T_993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1610;
  reg [31:0] _T_993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1611;
  reg [31:0] _T_994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1612;
  reg [31:0] _T_994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1613;
  reg [31:0] _T_995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1614;
  reg [31:0] _T_995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1615;
  reg [31:0] _T_996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1616;
  reg [31:0] _T_996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1617;
  reg [31:0] _T_997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1618;
  reg [31:0] _T_997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1619;
  reg [31:0] _T_998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1620;
  reg [31:0] _T_998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1621;
  reg [31:0] _T_999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1622;
  reg [31:0] _T_999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1623;
  reg [31:0] _T_1000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1624;
  reg [31:0] _T_1000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1625;
  reg [31:0] _T_1001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1626;
  reg [31:0] _T_1001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1627;
  reg [31:0] _T_1002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1628;
  reg [31:0] _T_1002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1629;
  reg [31:0] _T_1003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1630;
  reg [31:0] _T_1003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1631;
  reg [31:0] _T_1004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1632;
  reg [31:0] _T_1004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1633;
  reg [31:0] _T_1005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1634;
  reg [31:0] _T_1005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1635;
  reg [31:0] _T_1006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1636;
  reg [31:0] _T_1006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1637;
  reg [31:0] _T_1007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1638;
  reg [31:0] _T_1007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1639;
  reg [31:0] _T_1008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1640;
  reg [31:0] _T_1008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1641;
  reg [31:0] _T_1009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1642;
  reg [31:0] _T_1009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1643;
  reg [31:0] _T_1010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1644;
  reg [31:0] _T_1010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1645;
  reg [31:0] _T_1011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1646;
  reg [31:0] _T_1011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1647;
  reg [31:0] _T_1012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1648;
  reg [31:0] _T_1012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1649;
  reg [31:0] _T_1013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1650;
  reg [31:0] _T_1013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1651;
  reg [31:0] _T_1014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1652;
  reg [31:0] _T_1014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1653;
  reg [31:0] _T_1015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1654;
  reg [31:0] _T_1015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1655;
  reg [31:0] _T_1016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1656;
  reg [31:0] _T_1016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1657;
  reg [31:0] _T_1017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1658;
  reg [31:0] _T_1017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1659;
  reg [31:0] _T_1018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1660;
  reg [31:0] _T_1018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1661;
  reg [31:0] _T_1019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1662;
  reg [31:0] _T_1019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1663;
  reg [31:0] _T_1020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1664;
  reg [31:0] _T_1020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1665;
  reg [31:0] _T_1021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1666;
  reg [31:0] _T_1021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1667;
  reg [31:0] _T_1022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1668;
  reg [31:0] _T_1022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1669;
  reg [31:0] _T_1023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1670;
  reg [31:0] _T_1023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1671;
  reg [31:0] _T_1024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1672;
  reg [31:0] _T_1024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1673;
  reg [31:0] _T_1025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1674;
  reg [31:0] _T_1025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1675;
  reg [31:0] _T_1026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1676;
  reg [31:0] _T_1026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1677;
  reg [31:0] _T_1027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1678;
  reg [31:0] _T_1027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1679;
  reg [31:0] _T_1028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1680;
  reg [31:0] _T_1028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1681;
  reg [31:0] _T_1029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1682;
  reg [31:0] _T_1029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1683;
  reg [31:0] _T_1030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1684;
  reg [31:0] _T_1030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1685;
  reg [31:0] _T_1031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1686;
  reg [31:0] _T_1031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1687;
  reg [31:0] _T_1032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1688;
  reg [31:0] _T_1032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1689;
  reg [31:0] _T_1033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1690;
  reg [31:0] _T_1033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1691;
  reg [31:0] _T_1034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1692;
  reg [31:0] _T_1034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1693;
  reg [31:0] _T_1035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1694;
  reg [31:0] _T_1035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1695;
  reg [31:0] _T_1036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1696;
  reg [31:0] _T_1036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1697;
  reg [31:0] _T_1037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1698;
  reg [31:0] _T_1037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1699;
  reg [31:0] _T_1038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1700;
  reg [31:0] _T_1038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1701;
  reg [31:0] _T_1039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1702;
  reg [31:0] _T_1039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1703;
  reg [31:0] _T_1040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1704;
  reg [31:0] _T_1040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1705;
  reg [31:0] _T_1041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1706;
  reg [31:0] _T_1041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1707;
  reg [31:0] _T_1042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1708;
  reg [31:0] _T_1042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1709;
  reg [31:0] _T_1043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1710;
  reg [31:0] _T_1043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1711;
  reg [31:0] _T_1044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1712;
  reg [31:0] _T_1044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1713;
  reg [31:0] _T_1045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1714;
  reg [31:0] _T_1045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1715;
  reg [31:0] _T_1046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1716;
  reg [31:0] _T_1046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1717;
  reg [31:0] _T_1047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1718;
  reg [31:0] _T_1047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1719;
  reg [31:0] _T_1048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1720;
  reg [31:0] _T_1048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1721;
  reg [31:0] _T_1049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1722;
  reg [31:0] _T_1049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1723;
  reg [31:0] _T_1050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1724;
  reg [31:0] _T_1050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1725;
  reg [31:0] _T_1051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1726;
  reg [31:0] _T_1051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1727;
  reg [31:0] _T_1052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1728;
  reg [31:0] _T_1052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1729;
  reg [31:0] _T_1053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1730;
  reg [31:0] _T_1053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1731;
  reg [31:0] _T_1054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1732;
  reg [31:0] _T_1054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1733;
  reg [31:0] _T_1055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1734;
  reg [31:0] _T_1055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1735;
  reg [31:0] _T_1056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1736;
  reg [31:0] _T_1056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1737;
  reg [31:0] _T_1057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1738;
  reg [31:0] _T_1057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1739;
  reg [31:0] _T_1058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1740;
  reg [31:0] _T_1058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1741;
  reg [31:0] _T_1059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1742;
  reg [31:0] _T_1059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1743;
  reg [31:0] _T_1060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1744;
  reg [31:0] _T_1060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1745;
  reg [31:0] _T_1061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1746;
  reg [31:0] _T_1061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1747;
  reg [31:0] _T_1062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1748;
  reg [31:0] _T_1062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1749;
  reg [31:0] _T_1063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1750;
  reg [31:0] _T_1063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1751;
  reg [31:0] _T_1064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1752;
  reg [31:0] _T_1064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1753;
  reg [31:0] _T_1065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1754;
  reg [31:0] _T_1065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1755;
  reg [31:0] _T_1066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1756;
  reg [31:0] _T_1066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1757;
  reg [31:0] _T_1067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1758;
  reg [31:0] _T_1067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1759;
  reg [31:0] _T_1068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1760;
  reg [31:0] _T_1068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1761;
  reg [31:0] _T_1069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1762;
  reg [31:0] _T_1069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1763;
  reg [31:0] _T_1070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1764;
  reg [31:0] _T_1070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1765;
  reg [31:0] _T_1071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1766;
  reg [31:0] _T_1071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1767;
  reg [31:0] _T_1072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1768;
  reg [31:0] _T_1072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1769;
  reg [31:0] _T_1073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1770;
  reg [31:0] _T_1073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1771;
  reg [31:0] _T_1074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1772;
  reg [31:0] _T_1074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1773;
  reg [31:0] _T_1075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1774;
  reg [31:0] _T_1075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1775;
  reg [31:0] _T_1076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1776;
  reg [31:0] _T_1076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1777;
  reg [31:0] _T_1077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1778;
  reg [31:0] _T_1077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1779;
  reg [31:0] _T_1078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1780;
  reg [31:0] _T_1078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1781;
  reg [31:0] _T_1079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1782;
  reg [31:0] _T_1079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1783;
  reg [31:0] _T_1080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1784;
  reg [31:0] _T_1080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1785;
  reg [31:0] _T_1081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1786;
  reg [31:0] _T_1081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1787;
  reg [31:0] _T_1082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1788;
  reg [31:0] _T_1082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1789;
  reg [31:0] _T_1083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1790;
  reg [31:0] _T_1083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1791;
  reg [31:0] _T_1084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1792;
  reg [31:0] _T_1084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1793;
  reg [31:0] _T_1085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1794;
  reg [31:0] _T_1085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1795;
  reg [31:0] _T_1086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1796;
  reg [31:0] _T_1086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1797;
  reg [31:0] _T_1087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1798;
  reg [31:0] _T_1087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1799;
  reg [31:0] _T_1088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1800;
  reg [31:0] _T_1088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1801;
  reg [31:0] _T_1089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1802;
  reg [31:0] _T_1089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1803;
  reg [31:0] _T_1090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1804;
  reg [31:0] _T_1090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1805;
  reg [31:0] _T_1091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1806;
  reg [31:0] _T_1091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1807;
  reg [31:0] _T_1092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1808;
  reg [31:0] _T_1092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1809;
  reg [31:0] _T_1093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1810;
  reg [31:0] _T_1093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1811;
  reg [31:0] _T_1094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1812;
  reg [31:0] _T_1094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1813;
  reg [31:0] _T_1095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1814;
  reg [31:0] _T_1095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1815;
  reg [31:0] _T_1096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1816;
  reg [31:0] _T_1096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1817;
  reg [31:0] _T_1097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1818;
  reg [31:0] _T_1097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1819;
  reg [31:0] _T_1098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1820;
  reg [31:0] _T_1098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1821;
  reg [31:0] _T_1099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1822;
  reg [31:0] _T_1099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1823;
  reg [31:0] _T_1100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1824;
  reg [31:0] _T_1100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1825;
  reg [31:0] _T_1101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1826;
  reg [31:0] _T_1101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1827;
  reg [31:0] _T_1102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1828;
  reg [31:0] _T_1102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1829;
  reg [31:0] _T_1103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1830;
  reg [31:0] _T_1103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1831;
  reg [31:0] _T_1104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1832;
  reg [31:0] _T_1104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1833;
  reg [31:0] _T_1105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1834;
  reg [31:0] _T_1105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1835;
  reg [31:0] _T_1106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1836;
  reg [31:0] _T_1106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1837;
  reg [31:0] _T_1107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1838;
  reg [31:0] _T_1107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1839;
  reg [31:0] _T_1108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1840;
  reg [31:0] _T_1108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1841;
  reg [31:0] _T_1109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1842;
  reg [31:0] _T_1109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1843;
  reg [31:0] _T_1110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1844;
  reg [31:0] _T_1110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1845;
  reg [31:0] _T_1111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1846;
  reg [31:0] _T_1111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1847;
  reg [31:0] _T_1112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1848;
  reg [31:0] _T_1112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1849;
  reg [31:0] _T_1113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1850;
  reg [31:0] _T_1113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1851;
  reg [31:0] _T_1114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1852;
  reg [31:0] _T_1114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1853;
  reg [31:0] _T_1115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1854;
  reg [31:0] _T_1115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1855;
  reg [31:0] _T_1116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1856;
  reg [31:0] _T_1116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1857;
  reg [31:0] _T_1117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1858;
  reg [31:0] _T_1117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1859;
  reg [31:0] _T_1118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1860;
  reg [31:0] _T_1118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1861;
  reg [31:0] _T_1119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1862;
  reg [31:0] _T_1119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1863;
  reg [31:0] _T_1120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1864;
  reg [31:0] _T_1120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1865;
  reg [31:0] _T_1121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1866;
  reg [31:0] _T_1121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1867;
  reg [31:0] _T_1122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1868;
  reg [31:0] _T_1122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1869;
  reg [31:0] _T_1123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1870;
  reg [31:0] _T_1123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1871;
  reg [31:0] _T_1124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1872;
  reg [31:0] _T_1124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1873;
  reg [31:0] _T_1125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1874;
  reg [31:0] _T_1125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1875;
  reg [31:0] _T_1126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1876;
  reg [31:0] _T_1126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1877;
  reg [31:0] _T_1127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1878;
  reg [31:0] _T_1127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1879;
  reg [31:0] _T_1128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1880;
  reg [31:0] _T_1128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1881;
  reg [31:0] _T_1129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1882;
  reg [31:0] _T_1129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1883;
  reg [31:0] _T_1130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1884;
  reg [31:0] _T_1130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1885;
  reg [31:0] _T_1131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1886;
  reg [31:0] _T_1131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1887;
  reg [31:0] _T_1132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1888;
  reg [31:0] _T_1132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1889;
  reg [31:0] _T_1133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1890;
  reg [31:0] _T_1133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1891;
  reg [31:0] _T_1134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1892;
  reg [31:0] _T_1134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1893;
  reg [31:0] _T_1135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1894;
  reg [31:0] _T_1135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1895;
  reg [31:0] _T_1136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1896;
  reg [31:0] _T_1136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1897;
  reg [31:0] _T_1137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1898;
  reg [31:0] _T_1137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1899;
  reg [31:0] _T_1138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1900;
  reg [31:0] _T_1138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1901;
  reg [31:0] _T_1139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1902;
  reg [31:0] _T_1139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1903;
  reg [31:0] _T_1140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1904;
  reg [31:0] _T_1140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1905;
  reg [31:0] _T_1141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1906;
  reg [31:0] _T_1141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1907;
  reg [31:0] _T_1142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1908;
  reg [31:0] _T_1142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1909;
  reg [31:0] _T_1143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1910;
  reg [31:0] _T_1143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1911;
  reg [31:0] _T_1144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1912;
  reg [31:0] _T_1144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1913;
  reg [31:0] _T_1145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1914;
  reg [31:0] _T_1145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1915;
  reg [31:0] _T_1146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1916;
  reg [31:0] _T_1146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1917;
  reg [31:0] _T_1147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1918;
  reg [31:0] _T_1147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1919;
  reg [31:0] _T_1148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1920;
  reg [31:0] _T_1148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1921;
  reg [31:0] _T_1149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1922;
  reg [31:0] _T_1149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1923;
  reg [31:0] _T_1150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1924;
  reg [31:0] _T_1150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1925;
  reg [31:0] _T_1151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1926;
  reg [31:0] _T_1151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1927;
  reg [31:0] _T_1152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1928;
  reg [31:0] _T_1152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1929;
  reg [31:0] _T_1153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1930;
  reg [31:0] _T_1153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1931;
  reg [31:0] _T_1154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1932;
  reg [31:0] _T_1154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1933;
  reg [31:0] _T_1155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1934;
  reg [31:0] _T_1155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1935;
  reg [31:0] _T_1156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1936;
  reg [31:0] _T_1156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1937;
  reg [31:0] _T_1157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1938;
  reg [31:0] _T_1157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1939;
  reg [31:0] _T_1158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1940;
  reg [31:0] _T_1158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1941;
  reg [31:0] _T_1159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1942;
  reg [31:0] _T_1159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1943;
  reg [31:0] _T_1160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1944;
  reg [31:0] _T_1160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1945;
  reg [31:0] _T_1161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1946;
  reg [31:0] _T_1161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1947;
  reg [31:0] _T_1162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1948;
  reg [31:0] _T_1162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1949;
  reg [31:0] _T_1163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1950;
  reg [31:0] _T_1163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1951;
  reg [31:0] _T_1164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1952;
  reg [31:0] _T_1164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1953;
  reg [31:0] _T_1165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1954;
  reg [31:0] _T_1165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1955;
  reg [31:0] _T_1166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1956;
  reg [31:0] _T_1166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1957;
  reg [31:0] _T_1167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1958;
  reg [31:0] _T_1167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1959;
  reg [31:0] _T_1168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1960;
  reg [31:0] _T_1168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1961;
  reg [31:0] _T_1169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1962;
  reg [31:0] _T_1169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1963;
  reg [31:0] _T_1170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1964;
  reg [31:0] _T_1170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1965;
  reg [31:0] _T_1171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1966;
  reg [31:0] _T_1171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1967;
  reg [31:0] _T_1172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1968;
  reg [31:0] _T_1172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1969;
  reg [31:0] _T_1173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1970;
  reg [31:0] _T_1173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1971;
  reg [31:0] _T_1174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1972;
  reg [31:0] _T_1174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1973;
  reg [31:0] _T_1175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1974;
  reg [31:0] _T_1175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1975;
  reg [31:0] _T_1176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1976;
  reg [31:0] _T_1176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1977;
  reg [31:0] _T_1177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1978;
  reg [31:0] _T_1177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1979;
  reg [31:0] _T_1178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1980;
  reg [31:0] _T_1178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1981;
  reg [31:0] _T_1179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1982;
  reg [31:0] _T_1179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1983;
  reg [31:0] _T_1180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1984;
  reg [31:0] _T_1180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1985;
  reg [31:0] _T_1181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1986;
  reg [31:0] _T_1181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1987;
  reg [31:0] _T_1182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1988;
  reg [31:0] _T_1182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1989;
  reg [31:0] _T_1183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1990;
  reg [31:0] _T_1183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1991;
  reg [31:0] _T_1184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1992;
  reg [31:0] _T_1184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1993;
  reg [31:0] _T_1185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1994;
  reg [31:0] _T_1185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1995;
  reg [31:0] _T_1186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1996;
  reg [31:0] _T_1186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1997;
  reg [31:0] _T_1187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1998;
  reg [31:0] _T_1187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1999;
  reg [31:0] _T_1188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2000;
  reg [31:0] _T_1188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2001;
  reg [31:0] _T_1189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2002;
  reg [31:0] _T_1189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2003;
  reg [31:0] _T_1190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2004;
  reg [31:0] _T_1190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2005;
  reg [31:0] _T_1191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2006;
  reg [31:0] _T_1191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2007;
  reg [31:0] _T_1192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2008;
  reg [31:0] _T_1192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2009;
  reg [31:0] _T_1193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2010;
  reg [31:0] _T_1193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2011;
  reg [31:0] _T_1194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2012;
  reg [31:0] _T_1194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2013;
  reg [31:0] _T_1195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2014;
  reg [31:0] _T_1195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2015;
  reg [31:0] _T_1196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2016;
  reg [31:0] _T_1196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2017;
  reg [31:0] _T_1197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2018;
  reg [31:0] _T_1197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2019;
  reg [31:0] _T_1198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2020;
  reg [31:0] _T_1198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2021;
  reg [31:0] _T_1199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2022;
  reg [31:0] _T_1199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2023;
  reg [31:0] _T_1200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2024;
  reg [31:0] _T_1200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2025;
  reg [31:0] _T_1201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2026;
  reg [31:0] _T_1201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2027;
  reg [31:0] _T_1202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2028;
  reg [31:0] _T_1202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2029;
  reg [31:0] _T_1203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2030;
  reg [31:0] _T_1203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2031;
  reg [31:0] _T_1204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2032;
  reg [31:0] _T_1204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2033;
  reg [31:0] _T_1205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2034;
  reg [31:0] _T_1205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2035;
  reg [31:0] _T_1206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2036;
  reg [31:0] _T_1206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2037;
  reg [31:0] _T_1207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2038;
  reg [31:0] _T_1207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2039;
  reg [31:0] _T_1208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2040;
  reg [31:0] _T_1208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2041;
  reg [31:0] _T_1209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2042;
  reg [31:0] _T_1209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2043;
  reg [31:0] _T_1210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2044;
  reg [31:0] _T_1210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2045;
  reg [31:0] _T_1211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2046;
  reg [31:0] _T_1211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2047;
  reg [31:0] _T_1212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2048;
  reg [31:0] _T_1212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2049;
  reg [31:0] _T_1213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2050;
  reg [31:0] _T_1213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2051;
  reg [31:0] _T_1214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2052;
  reg [31:0] _T_1214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2053;
  reg [31:0] _T_1215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2054;
  reg [31:0] _T_1215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2055;
  reg [31:0] _T_1216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2056;
  reg [31:0] _T_1216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2057;
  reg [31:0] _T_1217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2058;
  reg [31:0] _T_1217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2059;
  reg [31:0] _T_1218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2060;
  reg [31:0] _T_1218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2061;
  reg [31:0] _T_1219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2062;
  reg [31:0] _T_1219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2063;
  reg [31:0] _T_1220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2064;
  reg [31:0] _T_1220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2065;
  reg [31:0] _T_1221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2066;
  reg [31:0] _T_1221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2067;
  reg [31:0] _T_1222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2068;
  reg [31:0] _T_1222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2069;
  reg [31:0] _T_1223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2070;
  reg [31:0] _T_1223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2071;
  reg [31:0] _T_1224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2072;
  reg [31:0] _T_1224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2073;
  reg [31:0] _T_1225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2074;
  reg [31:0] _T_1225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2075;
  reg [31:0] _T_1226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2076;
  reg [31:0] _T_1226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2077;
  reg [31:0] _T_1227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2078;
  reg [31:0] _T_1227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2079;
  reg [31:0] _T_1228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2080;
  reg [31:0] _T_1228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2081;
  reg [31:0] _T_1229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2082;
  reg [31:0] _T_1229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2083;
  reg [31:0] _T_1230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2084;
  reg [31:0] _T_1230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2085;
  reg [31:0] _T_1231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2086;
  reg [31:0] _T_1231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2087;
  reg [31:0] _T_1232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2088;
  reg [31:0] _T_1232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2089;
  reg [31:0] _T_1233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2090;
  reg [31:0] _T_1233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2091;
  reg [31:0] _T_1234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2092;
  reg [31:0] _T_1234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2093;
  reg [31:0] _T_1235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2094;
  reg [31:0] _T_1235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2095;
  reg [31:0] _T_1236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2096;
  reg [31:0] _T_1236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2097;
  reg [31:0] _T_1237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2098;
  reg [31:0] _T_1237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2099;
  reg [31:0] _T_1238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2100;
  reg [31:0] _T_1238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2101;
  reg [31:0] _T_1239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2102;
  reg [31:0] _T_1239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2103;
  reg [31:0] _T_1240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2104;
  reg [31:0] _T_1240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2105;
  reg [31:0] _T_1241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2106;
  reg [31:0] _T_1241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2107;
  reg [31:0] _T_1242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2108;
  reg [31:0] _T_1242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2109;
  reg [31:0] _T_1243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2110;
  reg [31:0] _T_1243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2111;
  reg [31:0] _T_1244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2112;
  reg [31:0] _T_1244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2113;
  reg [31:0] _T_1245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2114;
  reg [31:0] _T_1245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2115;
  reg [31:0] _T_1246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2116;
  reg [31:0] _T_1246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2117;
  reg [31:0] _T_1247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2118;
  reg [31:0] _T_1247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2119;
  reg [31:0] _T_1248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2120;
  reg [31:0] _T_1248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2121;
  reg [31:0] _T_1249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2122;
  reg [31:0] _T_1249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2123;
  reg [31:0] _T_1250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2124;
  reg [31:0] _T_1250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2125;
  reg [31:0] _T_1251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2126;
  reg [31:0] _T_1251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2127;
  reg [31:0] _T_1252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2128;
  reg [31:0] _T_1252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2129;
  reg [31:0] _T_1253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2130;
  reg [31:0] _T_1253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2131;
  reg [31:0] _T_1254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2132;
  reg [31:0] _T_1254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2133;
  reg [31:0] _T_1255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2134;
  reg [31:0] _T_1255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2135;
  reg [31:0] _T_1256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2136;
  reg [31:0] _T_1256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2137;
  reg [31:0] _T_1257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2138;
  reg [31:0] _T_1257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2139;
  reg [31:0] _T_1258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2140;
  reg [31:0] _T_1258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2141;
  reg [31:0] _T_1259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2142;
  reg [31:0] _T_1259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2143;
  reg [31:0] _T_1260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2144;
  reg [31:0] _T_1260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2145;
  reg [31:0] _T_1261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2146;
  reg [31:0] _T_1261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2147;
  reg [31:0] _T_1262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2148;
  reg [31:0] _T_1262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2149;
  reg [31:0] _T_1263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2150;
  reg [31:0] _T_1263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2151;
  reg [31:0] _T_1264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2152;
  reg [31:0] _T_1264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2153;
  reg [31:0] _T_1265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2154;
  reg [31:0] _T_1265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2155;
  reg [31:0] _T_1266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2156;
  reg [31:0] _T_1266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2157;
  reg [31:0] _T_1267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2158;
  reg [31:0] _T_1267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2159;
  reg [31:0] _T_1268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2160;
  reg [31:0] _T_1268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2161;
  reg [31:0] _T_1269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2162;
  reg [31:0] _T_1269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2163;
  reg [31:0] _T_1270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2164;
  reg [31:0] _T_1270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2165;
  reg [31:0] _T_1271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2166;
  reg [31:0] _T_1271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2167;
  reg [31:0] _T_1272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2168;
  reg [31:0] _T_1272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2169;
  reg [31:0] _T_1273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2170;
  reg [31:0] _T_1273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2171;
  reg [31:0] _T_1274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2172;
  reg [31:0] _T_1274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2173;
  reg [31:0] _T_1275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2174;
  reg [31:0] _T_1275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2175;
  reg [31:0] _T_1276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2176;
  reg [31:0] _T_1276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2177;
  reg [31:0] _T_1277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2178;
  reg [31:0] _T_1277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2179;
  reg [31:0] _T_1278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2180;
  reg [31:0] _T_1278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2181;
  reg [31:0] _T_1279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2182;
  reg [31:0] _T_1279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2183;
  reg [31:0] _T_1280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2184;
  reg [31:0] _T_1280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2185;
  reg [31:0] _T_1281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2186;
  reg [31:0] _T_1281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2187;
  reg [31:0] _T_1282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2188;
  reg [31:0] _T_1282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2189;
  reg [31:0] _T_1283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2190;
  reg [31:0] _T_1283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2191;
  reg [31:0] _T_1284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2192;
  reg [31:0] _T_1284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2193;
  reg [31:0] _T_1285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2194;
  reg [31:0] _T_1285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2195;
  reg [31:0] _T_1286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2196;
  reg [31:0] _T_1286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2197;
  reg [31:0] _T_1287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2198;
  reg [31:0] _T_1287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2199;
  reg [31:0] _T_1288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2200;
  reg [31:0] _T_1288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2201;
  reg [31:0] _T_1289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2202;
  reg [31:0] _T_1289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2203;
  reg [31:0] _T_1290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2204;
  reg [31:0] _T_1290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2205;
  reg [31:0] _T_1291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2206;
  reg [31:0] _T_1291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2207;
  reg [31:0] _T_1292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2208;
  reg [31:0] _T_1292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2209;
  reg [31:0] _T_1293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2210;
  reg [31:0] _T_1293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2211;
  reg [31:0] _T_1294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2212;
  reg [31:0] _T_1294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2213;
  reg [31:0] _T_1295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2214;
  reg [31:0] _T_1295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2215;
  reg [31:0] _T_1296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2216;
  reg [31:0] _T_1296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2217;
  reg [31:0] _T_1297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2218;
  reg [31:0] _T_1297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2219;
  reg [31:0] _T_1298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2220;
  reg [31:0] _T_1298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2221;
  reg [31:0] _T_1299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2222;
  reg [31:0] _T_1299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2223;
  reg [31:0] _T_1300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2224;
  reg [31:0] _T_1300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2225;
  reg [31:0] _T_1301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2226;
  reg [31:0] _T_1301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2227;
  reg [31:0] _T_1302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2228;
  reg [31:0] _T_1302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2229;
  reg [31:0] _T_1303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2230;
  reg [31:0] _T_1303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2231;
  reg [31:0] _T_1304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2232;
  reg [31:0] _T_1304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2233;
  reg [31:0] _T_1305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2234;
  reg [31:0] _T_1305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2235;
  reg [31:0] _T_1306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2236;
  reg [31:0] _T_1306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2237;
  reg [31:0] _T_1307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2238;
  reg [31:0] _T_1307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2239;
  reg [31:0] _T_1308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2240;
  reg [31:0] _T_1308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2241;
  reg [31:0] _T_1309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2242;
  reg [31:0] _T_1309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2243;
  reg [31:0] _T_1310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2244;
  reg [31:0] _T_1310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2245;
  reg [31:0] _T_1311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2246;
  reg [31:0] _T_1311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2247;
  reg [31:0] _T_1312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2248;
  reg [31:0] _T_1312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2249;
  reg [31:0] _T_1313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2250;
  reg [31:0] _T_1313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2251;
  reg [31:0] _T_1314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2252;
  reg [31:0] _T_1314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2253;
  reg [31:0] _T_1315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2254;
  reg [31:0] _T_1315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2255;
  reg [31:0] _T_1316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2256;
  reg [31:0] _T_1316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2257;
  reg [31:0] _T_1317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2258;
  reg [31:0] _T_1317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2259;
  reg [31:0] _T_1318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2260;
  reg [31:0] _T_1318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2261;
  reg [31:0] _T_1319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2262;
  reg [31:0] _T_1319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2263;
  reg [31:0] _T_1320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2264;
  reg [31:0] _T_1320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2265;
  reg [31:0] _T_1321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2266;
  reg [31:0] _T_1321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2267;
  reg [31:0] _T_1322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2268;
  reg [31:0] _T_1322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2269;
  reg [31:0] _T_1323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2270;
  reg [31:0] _T_1323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2271;
  reg [31:0] _T_1324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2272;
  reg [31:0] _T_1324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2273;
  reg [31:0] _T_1325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2274;
  reg [31:0] _T_1325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2275;
  reg [31:0] _T_1326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2276;
  reg [31:0] _T_1326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2277;
  reg [31:0] _T_1327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2278;
  reg [31:0] _T_1327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2279;
  reg [31:0] _T_1328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2280;
  reg [31:0] _T_1328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2281;
  reg [31:0] _T_1329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2282;
  reg [31:0] _T_1329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2283;
  reg [31:0] _T_1330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2284;
  reg [31:0] _T_1330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2285;
  reg [31:0] _T_1331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2286;
  reg [31:0] _T_1331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2287;
  reg [31:0] _T_1332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2288;
  reg [31:0] _T_1332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2289;
  reg [31:0] _T_1333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2290;
  reg [31:0] _T_1333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2291;
  reg [31:0] _T_1334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2292;
  reg [31:0] _T_1334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2293;
  reg [31:0] _T_1335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2294;
  reg [31:0] _T_1335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2295;
  reg [31:0] _T_1336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2296;
  reg [31:0] _T_1336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2297;
  reg [31:0] _T_1337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2298;
  reg [31:0] _T_1337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2299;
  reg [31:0] _T_1338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2300;
  reg [31:0] _T_1338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2301;
  reg [31:0] _T_1339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2302;
  reg [31:0] _T_1339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2303;
  reg [31:0] _T_1340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2304;
  reg [31:0] _T_1340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2305;
  reg [31:0] _T_1341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2306;
  reg [31:0] _T_1341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2307;
  reg [31:0] _T_1342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2308;
  reg [31:0] _T_1342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2309;
  reg [31:0] _T_1343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2310;
  reg [31:0] _T_1343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2311;
  reg [31:0] _T_1344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2312;
  reg [31:0] _T_1344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2313;
  reg [31:0] _T_1345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2314;
  reg [31:0] _T_1345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2315;
  reg [31:0] _T_1346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2316;
  reg [31:0] _T_1346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2317;
  reg [31:0] _T_1347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2318;
  reg [31:0] _T_1347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2319;
  reg [31:0] _T_1348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2320;
  reg [31:0] _T_1348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2321;
  reg [31:0] _T_1349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2322;
  reg [31:0] _T_1349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2323;
  reg [31:0] _T_1350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2324;
  reg [31:0] _T_1350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2325;
  reg [31:0] _T_1351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2326;
  reg [31:0] _T_1351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2327;
  reg [31:0] _T_1352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2328;
  reg [31:0] _T_1352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2329;
  reg [31:0] _T_1353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2330;
  reg [31:0] _T_1353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2331;
  reg [31:0] _T_1354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2332;
  reg [31:0] _T_1354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2333;
  reg [31:0] _T_1355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2334;
  reg [31:0] _T_1355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2335;
  reg [31:0] _T_1356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2336;
  reg [31:0] _T_1356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2337;
  reg [31:0] _T_1357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2338;
  reg [31:0] _T_1357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2339;
  reg [31:0] _T_1358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2340;
  reg [31:0] _T_1358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2341;
  reg [31:0] _T_1359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2342;
  reg [31:0] _T_1359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2343;
  reg [31:0] _T_1360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2344;
  reg [31:0] _T_1360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2345;
  reg [31:0] _T_1361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2346;
  reg [31:0] _T_1361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2347;
  reg [31:0] _T_1362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2348;
  reg [31:0] _T_1362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2349;
  reg [31:0] _T_1363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2350;
  reg [31:0] _T_1363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2351;
  reg [31:0] _T_1364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2352;
  reg [31:0] _T_1364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2353;
  reg [31:0] _T_1365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2354;
  reg [31:0] _T_1365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2355;
  reg [31:0] _T_1366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2356;
  reg [31:0] _T_1366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2357;
  reg [31:0] _T_1367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2358;
  reg [31:0] _T_1367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2359;
  reg [31:0] _T_1368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2360;
  reg [31:0] _T_1368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2361;
  reg [31:0] _T_1369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2362;
  reg [31:0] _T_1369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2363;
  reg [31:0] _T_1370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2364;
  reg [31:0] _T_1370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2365;
  reg [31:0] _T_1371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2366;
  reg [31:0] _T_1371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2367;
  reg [31:0] _T_1372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2368;
  reg [31:0] _T_1372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2369;
  reg [31:0] _T_1373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2370;
  reg [31:0] _T_1373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2371;
  reg [31:0] _T_1374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2372;
  reg [31:0] _T_1374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2373;
  reg [31:0] _T_1375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2374;
  reg [31:0] _T_1375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2375;
  reg [31:0] _T_1376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2376;
  reg [31:0] _T_1376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2377;
  reg [31:0] _T_1377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2378;
  reg [31:0] _T_1377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2379;
  reg [31:0] _T_1378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2380;
  reg [31:0] _T_1378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2381;
  reg [31:0] _T_1379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2382;
  reg [31:0] _T_1379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2383;
  reg [31:0] _T_1380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2384;
  reg [31:0] _T_1380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2385;
  reg [31:0] _T_1381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2386;
  reg [31:0] _T_1381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2387;
  reg [31:0] _T_1382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2388;
  reg [31:0] _T_1382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2389;
  reg [31:0] _T_1383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2390;
  reg [31:0] _T_1383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2391;
  reg [31:0] _T_1384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2392;
  reg [31:0] _T_1384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2393;
  reg [31:0] _T_1385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2394;
  reg [31:0] _T_1385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2395;
  reg [31:0] _T_1386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2396;
  reg [31:0] _T_1386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2397;
  reg [31:0] _T_1387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2398;
  reg [31:0] _T_1387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2399;
  reg [31:0] _T_1388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2400;
  reg [31:0] _T_1388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2401;
  reg [31:0] _T_1389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2402;
  reg [31:0] _T_1389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2403;
  reg [31:0] _T_1390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2404;
  reg [31:0] _T_1390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2405;
  reg [31:0] _T_1391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2406;
  reg [31:0] _T_1391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2407;
  reg [31:0] _T_1392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2408;
  reg [31:0] _T_1392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2409;
  reg [31:0] _T_1393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2410;
  reg [31:0] _T_1393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2411;
  reg [31:0] _T_1394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2412;
  reg [31:0] _T_1394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2413;
  reg [31:0] _T_1395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2414;
  reg [31:0] _T_1395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2415;
  reg [31:0] _T_1396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2416;
  reg [31:0] _T_1396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2417;
  reg [31:0] _T_1397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2418;
  reg [31:0] _T_1397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2419;
  reg [31:0] _T_1398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2420;
  reg [31:0] _T_1398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2421;
  reg [31:0] _T_1399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2422;
  reg [31:0] _T_1399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2423;
  reg [31:0] _T_1400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2424;
  reg [31:0] _T_1400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2425;
  reg [31:0] _T_1401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2426;
  reg [31:0] _T_1401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2427;
  reg [31:0] _T_1402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2428;
  reg [31:0] _T_1402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2429;
  reg [31:0] _T_1403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2430;
  reg [31:0] _T_1403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2431;
  reg [31:0] _T_1404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2432;
  reg [31:0] _T_1404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2433;
  reg [31:0] _T_1405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2434;
  reg [31:0] _T_1405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2435;
  reg [31:0] _T_1406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2436;
  reg [31:0] _T_1406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2437;
  reg [31:0] _T_1407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2438;
  reg [31:0] _T_1407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2439;
  reg [31:0] _T_1408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2440;
  reg [31:0] _T_1408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2441;
  reg [31:0] _T_1409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2442;
  reg [31:0] _T_1409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2443;
  reg [31:0] _T_1410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2444;
  reg [31:0] _T_1410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2445;
  reg [31:0] _T_1411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2446;
  reg [31:0] _T_1411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2447;
  reg [31:0] _T_1412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2448;
  reg [31:0] _T_1412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2449;
  reg [31:0] _T_1413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2450;
  reg [31:0] _T_1413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2451;
  reg [31:0] _T_1414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2452;
  reg [31:0] _T_1414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2453;
  reg [31:0] _T_1415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2454;
  reg [31:0] _T_1415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2455;
  reg [31:0] _T_1416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2456;
  reg [31:0] _T_1416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2457;
  reg [31:0] _T_1417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2458;
  reg [31:0] _T_1417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2459;
  reg [31:0] _T_1418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2460;
  reg [31:0] _T_1418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2461;
  reg [31:0] _T_1419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2462;
  reg [31:0] _T_1419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2463;
  reg [31:0] _T_1420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2464;
  reg [31:0] _T_1420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2465;
  reg [31:0] _T_1421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2466;
  reg [31:0] _T_1421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2467;
  reg [31:0] _T_1422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2468;
  reg [31:0] _T_1422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2469;
  reg [31:0] _T_1423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2470;
  reg [31:0] _T_1423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2471;
  reg [31:0] _T_1424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2472;
  reg [31:0] _T_1424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2473;
  reg [31:0] _T_1425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2474;
  reg [31:0] _T_1425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2475;
  reg [31:0] _T_1426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2476;
  reg [31:0] _T_1426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2477;
  reg [31:0] _T_1427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2478;
  reg [31:0] _T_1427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2479;
  reg [31:0] _T_1428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2480;
  reg [31:0] _T_1428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2481;
  reg [31:0] _T_1429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2482;
  reg [31:0] _T_1429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2483;
  reg [31:0] _T_1430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2484;
  reg [31:0] _T_1430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2485;
  reg [31:0] _T_1431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2486;
  reg [31:0] _T_1431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2487;
  reg [31:0] _T_1432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2488;
  reg [31:0] _T_1432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2489;
  reg [31:0] _T_1433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2490;
  reg [31:0] _T_1433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2491;
  reg [31:0] _T_1434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2492;
  reg [31:0] _T_1434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2493;
  reg [31:0] _T_1435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2494;
  reg [31:0] _T_1435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2495;
  reg [31:0] _T_1436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2496;
  reg [31:0] _T_1436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2497;
  reg [31:0] _T_1437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2498;
  reg [31:0] _T_1437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2499;
  reg [31:0] _T_1438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2500;
  reg [31:0] _T_1438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2501;
  reg [31:0] _T_1439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2502;
  reg [31:0] _T_1439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2503;
  reg [31:0] _T_1440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2504;
  reg [31:0] _T_1440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2505;
  reg [31:0] _T_1441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2506;
  reg [31:0] _T_1441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2507;
  reg [31:0] _T_1442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2508;
  reg [31:0] _T_1442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2509;
  reg [31:0] _T_1443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2510;
  reg [31:0] _T_1443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2511;
  reg [31:0] _T_1444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2512;
  reg [31:0] _T_1444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2513;
  reg [31:0] _T_1445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2514;
  reg [31:0] _T_1445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2515;
  reg [31:0] _T_1446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2516;
  reg [31:0] _T_1446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2517;
  reg [31:0] _T_1447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2518;
  reg [31:0] _T_1447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2519;
  reg [31:0] _T_1448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2520;
  reg [31:0] _T_1448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2521;
  reg [31:0] _T_1449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2522;
  reg [31:0] _T_1449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2523;
  reg [31:0] _T_1450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2524;
  reg [31:0] _T_1450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2525;
  reg [31:0] _T_1451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2526;
  reg [31:0] _T_1451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2527;
  reg [31:0] _T_1452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2528;
  reg [31:0] _T_1452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2529;
  reg [31:0] _T_1453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2530;
  reg [31:0] _T_1453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2531;
  reg [31:0] _T_1454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2532;
  reg [31:0] _T_1454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2533;
  reg [31:0] _T_1455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2534;
  reg [31:0] _T_1455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2535;
  reg [31:0] _T_1456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2536;
  reg [31:0] _T_1456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2537;
  reg [31:0] _T_1457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2538;
  reg [31:0] _T_1457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2539;
  reg [31:0] _T_1458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2540;
  reg [31:0] _T_1458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2541;
  reg [31:0] _T_1459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2542;
  reg [31:0] _T_1459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2543;
  reg [31:0] _T_1460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2544;
  reg [31:0] _T_1460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2545;
  reg [31:0] _T_1461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2546;
  reg [31:0] _T_1461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2547;
  reg [31:0] _T_1462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2548;
  reg [31:0] _T_1462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2549;
  reg [31:0] _T_1463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2550;
  reg [31:0] _T_1463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2551;
  reg [31:0] _T_1464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2552;
  reg [31:0] _T_1464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2553;
  reg [31:0] _T_1465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2554;
  reg [31:0] _T_1465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2555;
  reg [31:0] _T_1466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2556;
  reg [31:0] _T_1466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2557;
  reg [31:0] _T_1467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2558;
  reg [31:0] _T_1467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2559;
  reg [31:0] _T_1468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2560;
  reg [31:0] _T_1468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2561;
  reg [31:0] _T_1469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2562;
  reg [31:0] _T_1469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2563;
  reg [31:0] _T_1470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2564;
  reg [31:0] _T_1470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2565;
  reg [31:0] _T_1471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2566;
  reg [31:0] _T_1471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2567;
  reg [31:0] _T_1472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2568;
  reg [31:0] _T_1472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2569;
  reg [31:0] _T_1473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2570;
  reg [31:0] _T_1473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2571;
  reg [31:0] _T_1474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2572;
  reg [31:0] _T_1474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2573;
  reg [31:0] _T_1475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2574;
  reg [31:0] _T_1475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2575;
  reg [31:0] _T_1476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2576;
  reg [31:0] _T_1476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2577;
  reg [31:0] _T_1477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2578;
  reg [31:0] _T_1477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2579;
  reg [31:0] _T_1478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2580;
  reg [31:0] _T_1478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2581;
  reg [31:0] _T_1479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2582;
  reg [31:0] _T_1479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2583;
  reg [31:0] _T_1480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2584;
  reg [31:0] _T_1480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2585;
  reg [31:0] _T_1481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2586;
  reg [31:0] _T_1481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2587;
  reg [31:0] _T_1482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2588;
  reg [31:0] _T_1482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2589;
  reg [31:0] _T_1483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2590;
  reg [31:0] _T_1483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2591;
  reg [31:0] _T_1484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2592;
  reg [31:0] _T_1484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2593;
  reg [31:0] _T_1485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2594;
  reg [31:0] _T_1485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2595;
  reg [31:0] _T_1486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2596;
  reg [31:0] _T_1486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2597;
  reg [31:0] _T_1487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2598;
  reg [31:0] _T_1487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2599;
  reg [31:0] _T_1488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2600;
  reg [31:0] _T_1488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2601;
  reg [31:0] _T_1489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2602;
  reg [31:0] _T_1489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2603;
  reg [31:0] _T_1490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2604;
  reg [31:0] _T_1490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2605;
  reg [31:0] _T_1491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2606;
  reg [31:0] _T_1491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2607;
  reg [31:0] _T_1492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2608;
  reg [31:0] _T_1492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2609;
  reg [31:0] _T_1493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2610;
  reg [31:0] _T_1493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2611;
  reg [31:0] _T_1494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2612;
  reg [31:0] _T_1494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2613;
  reg [31:0] _T_1495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2614;
  reg [31:0] _T_1495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2615;
  reg [31:0] _T_1496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2616;
  reg [31:0] _T_1496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2617;
  reg [31:0] _T_1497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2618;
  reg [31:0] _T_1497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2619;
  reg [31:0] _T_1498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2620;
  reg [31:0] _T_1498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2621;
  reg [31:0] _T_1499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2622;
  reg [31:0] _T_1499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2623;
  reg [31:0] _T_1500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2624;
  reg [31:0] _T_1500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2625;
  reg [31:0] _T_1501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2626;
  reg [31:0] _T_1501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2627;
  reg [31:0] _T_1502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2628;
  reg [31:0] _T_1502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2629;
  reg [31:0] _T_1503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2630;
  reg [31:0] _T_1503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2631;
  reg [31:0] _T_1504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2632;
  reg [31:0] _T_1504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2633;
  reg [31:0] _T_1505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2634;
  reg [31:0] _T_1505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2635;
  reg [31:0] _T_1506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2636;
  reg [31:0] _T_1506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2637;
  reg [31:0] _T_1507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2638;
  reg [31:0] _T_1507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2639;
  reg [31:0] _T_1508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2640;
  reg [31:0] _T_1508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2641;
  reg [31:0] _T_1509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2642;
  reg [31:0] _T_1509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2643;
  reg [31:0] _T_1510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2644;
  reg [31:0] _T_1510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2645;
  reg [31:0] _T_1511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2646;
  reg [31:0] _T_1511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2647;
  reg [31:0] _T_1512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2648;
  reg [31:0] _T_1512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2649;
  reg [31:0] _T_1513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2650;
  reg [31:0] _T_1513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2651;
  reg [31:0] _T_1514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2652;
  reg [31:0] _T_1514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2653;
  reg [31:0] _T_1515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2654;
  reg [31:0] _T_1515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2655;
  reg [31:0] _T_1516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2656;
  reg [31:0] _T_1516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2657;
  reg [31:0] _T_1517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2658;
  reg [31:0] _T_1517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2659;
  reg [31:0] _T_1518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2660;
  reg [31:0] _T_1518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2661;
  reg [31:0] _T_1519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2662;
  reg [31:0] _T_1519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2663;
  reg [31:0] _T_1520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2664;
  reg [31:0] _T_1520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2665;
  reg [31:0] _T_1521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2666;
  reg [31:0] _T_1521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2667;
  reg [31:0] _T_1522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2668;
  reg [31:0] _T_1522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2669;
  reg [31:0] _T_1523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2670;
  reg [31:0] _T_1523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2671;
  reg [31:0] _T_1524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2672;
  reg [31:0] _T_1524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2673;
  reg [31:0] _T_1525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2674;
  reg [31:0] _T_1525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2675;
  reg [31:0] _T_1526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2676;
  reg [31:0] _T_1526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2677;
  reg [31:0] _T_1527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2678;
  reg [31:0] _T_1527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2679;
  reg [31:0] _T_1528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2680;
  reg [31:0] _T_1528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2681;
  reg [31:0] _T_1529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2682;
  reg [31:0] _T_1529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2683;
  reg [31:0] _T_1530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2684;
  reg [31:0] _T_1530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2685;
  reg [31:0] _T_1531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2686;
  reg [31:0] _T_1531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2687;
  reg [31:0] _T_1532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2688;
  reg [31:0] _T_1532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2689;
  reg [31:0] _T_1533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2690;
  reg [31:0] _T_1533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2691;
  reg [31:0] _T_1534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2692;
  reg [31:0] _T_1534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2693;
  reg [31:0] _T_1535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2694;
  reg [31:0] _T_1535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2695;
  reg [31:0] _T_1536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2696;
  reg [31:0] _T_1536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2697;
  reg [31:0] _T_1537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2698;
  reg [31:0] _T_1537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2699;
  reg [31:0] _T_1538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2700;
  reg [31:0] _T_1538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2701;
  reg [31:0] _T_1539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2702;
  reg [31:0] _T_1539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2703;
  reg [31:0] _T_1540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2704;
  reg [31:0] _T_1540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2705;
  reg [31:0] _T_1541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2706;
  reg [31:0] _T_1541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2707;
  reg [31:0] _T_1542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2708;
  reg [31:0] _T_1542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2709;
  reg [31:0] _T_1543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2710;
  reg [31:0] _T_1543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2711;
  reg [31:0] _T_1544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2712;
  reg [31:0] _T_1544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2713;
  reg [31:0] _T_1545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2714;
  reg [31:0] _T_1545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2715;
  reg [31:0] _T_1546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2716;
  reg [31:0] _T_1546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2717;
  reg [31:0] _T_1547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2718;
  reg [31:0] _T_1547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2719;
  reg [31:0] _T_1548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2720;
  reg [31:0] _T_1548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2721;
  reg [31:0] _T_1549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2722;
  reg [31:0] _T_1549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2723;
  reg [31:0] _T_1550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2724;
  reg [31:0] _T_1550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2725;
  reg [31:0] _T_1551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2726;
  reg [31:0] _T_1551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2727;
  reg [31:0] _T_1552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2728;
  reg [31:0] _T_1552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2729;
  reg [31:0] _T_1553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2730;
  reg [31:0] _T_1553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2731;
  reg [31:0] _T_1554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2732;
  reg [31:0] _T_1554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2733;
  reg [31:0] _T_1555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2734;
  reg [31:0] _T_1555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2735;
  reg [31:0] _T_1556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2736;
  reg [31:0] _T_1556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2737;
  reg [31:0] _T_1557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2738;
  reg [31:0] _T_1557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2739;
  reg [31:0] _T_1558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2740;
  reg [31:0] _T_1558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2741;
  reg [31:0] _T_1559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2742;
  reg [31:0] _T_1559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2743;
  reg [31:0] _T_1560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2744;
  reg [31:0] _T_1560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2745;
  reg [31:0] _T_1561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2746;
  reg [31:0] _T_1561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2747;
  reg [31:0] _T_1562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2748;
  reg [31:0] _T_1562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2749;
  reg [31:0] _T_1563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2750;
  reg [31:0] _T_1563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2751;
  reg [31:0] _T_1564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2752;
  reg [31:0] _T_1564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2753;
  reg [31:0] _T_1565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2754;
  reg [31:0] _T_1565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2755;
  reg [31:0] _T_1566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2756;
  reg [31:0] _T_1566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2757;
  reg [31:0] _T_1567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2758;
  reg [31:0] _T_1567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2759;
  reg [31:0] _T_1568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2760;
  reg [31:0] _T_1568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2761;
  reg [31:0] _T_1569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2762;
  reg [31:0] _T_1569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2763;
  reg [31:0] _T_1570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2764;
  reg [31:0] _T_1570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2765;
  reg [31:0] _T_1571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2766;
  reg [31:0] _T_1571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2767;
  reg [31:0] _T_1572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2768;
  reg [31:0] _T_1572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2769;
  reg [31:0] _T_1573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2770;
  reg [31:0] _T_1573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2771;
  reg [31:0] _T_1574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2772;
  reg [31:0] _T_1574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2773;
  reg [31:0] _T_1575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2774;
  reg [31:0] _T_1575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2775;
  reg [31:0] _T_1576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2776;
  reg [31:0] _T_1576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2777;
  reg [31:0] _T_1577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2778;
  reg [31:0] _T_1577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2779;
  reg [31:0] _T_1578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2780;
  reg [31:0] _T_1578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2781;
  reg [31:0] _T_1579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2782;
  reg [31:0] _T_1579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2783;
  reg [31:0] _T_1580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2784;
  reg [31:0] _T_1580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2785;
  reg [31:0] _T_1581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2786;
  reg [31:0] _T_1581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2787;
  reg [31:0] _T_1582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2788;
  reg [31:0] _T_1582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2789;
  reg [31:0] _T_1583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2790;
  reg [31:0] _T_1583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2791;
  reg [31:0] _T_1584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2792;
  reg [31:0] _T_1584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2793;
  reg [31:0] _T_1585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2794;
  reg [31:0] _T_1585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2795;
  reg [31:0] _T_1586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2796;
  reg [31:0] _T_1586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2797;
  reg [31:0] _T_1587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2798;
  reg [31:0] _T_1587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2799;
  reg [31:0] _T_1588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2800;
  reg [31:0] _T_1588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2801;
  reg [31:0] _T_1589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2802;
  reg [31:0] _T_1589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2803;
  reg [31:0] _T_1590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2804;
  reg [31:0] _T_1590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2805;
  reg [31:0] _T_1591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2806;
  reg [31:0] _T_1591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2807;
  reg [31:0] _T_1592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2808;
  reg [31:0] _T_1592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2809;
  reg [31:0] _T_1593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2810;
  reg [31:0] _T_1593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2811;
  reg [31:0] _T_1594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2812;
  reg [31:0] _T_1594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2813;
  reg [31:0] _T_1595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2814;
  reg [31:0] _T_1595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2815;
  reg [31:0] _T_1596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2816;
  reg [31:0] _T_1596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2817;
  reg [31:0] _T_1597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2818;
  reg [31:0] _T_1597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2819;
  reg [31:0] _T_1598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2820;
  reg [31:0] _T_1598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2821;
  reg [31:0] _T_1599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2822;
  reg [31:0] _T_1599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2823;
  reg [31:0] _T_1600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2824;
  reg [31:0] _T_1600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2825;
  reg [31:0] _T_1601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2826;
  reg [31:0] _T_1601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2827;
  reg [31:0] _T_1602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2828;
  reg [31:0] _T_1602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2829;
  reg [31:0] _T_1603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2830;
  reg [31:0] _T_1603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2831;
  reg [31:0] _T_1604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2832;
  reg [31:0] _T_1604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2833;
  reg [31:0] _T_1605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2834;
  reg [31:0] _T_1605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2835;
  reg [31:0] _T_1606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2836;
  reg [31:0] _T_1606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2837;
  reg [31:0] _T_1607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2838;
  reg [31:0] _T_1607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2839;
  reg [31:0] _T_1608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2840;
  reg [31:0] _T_1608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2841;
  reg [31:0] _T_1609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2842;
  reg [31:0] _T_1609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2843;
  reg [31:0] _T_1610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2844;
  reg [31:0] _T_1610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2845;
  reg [31:0] _T_1611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2846;
  reg [31:0] _T_1611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2847;
  reg [31:0] _T_1612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2848;
  reg [31:0] _T_1612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2849;
  reg [31:0] _T_1613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2850;
  reg [31:0] _T_1613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2851;
  reg [31:0] _T_1614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2852;
  reg [31:0] _T_1614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2853;
  reg [31:0] _T_1615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2854;
  reg [31:0] _T_1615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2855;
  reg [31:0] _T_1616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2856;
  reg [31:0] _T_1616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2857;
  reg [31:0] _T_1617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2858;
  reg [31:0] _T_1617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2859;
  reg [31:0] _T_1618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2860;
  reg [31:0] _T_1618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2861;
  reg [31:0] _T_1619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2862;
  reg [31:0] _T_1619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2863;
  reg [31:0] _T_1620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2864;
  reg [31:0] _T_1620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2865;
  reg [31:0] _T_1621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2866;
  reg [31:0] _T_1621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2867;
  reg [31:0] _T_1622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2868;
  reg [31:0] _T_1622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2869;
  reg [31:0] _T_1623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2870;
  reg [31:0] _T_1623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2871;
  reg [31:0] _T_1624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2872;
  reg [31:0] _T_1624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2873;
  reg [31:0] _T_1625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2874;
  reg [31:0] _T_1625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2875;
  reg [31:0] _T_1626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2876;
  reg [31:0] _T_1626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2877;
  reg [31:0] _T_1627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2878;
  reg [31:0] _T_1627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2879;
  reg [31:0] _T_1628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2880;
  reg [31:0] _T_1628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2881;
  reg [31:0] _T_1629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2882;
  reg [31:0] _T_1629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2883;
  reg [31:0] _T_1630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2884;
  reg [31:0] _T_1630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2885;
  reg [31:0] _T_1631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2886;
  reg [31:0] _T_1631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2887;
  reg [31:0] _T_1632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2888;
  reg [31:0] _T_1632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2889;
  reg [31:0] _T_1633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2890;
  reg [31:0] _T_1633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2891;
  reg [31:0] _T_1634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2892;
  reg [31:0] _T_1634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2893;
  reg [31:0] _T_1635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2894;
  reg [31:0] _T_1635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2895;
  reg [31:0] _T_1636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2896;
  reg [31:0] _T_1636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2897;
  reg [31:0] _T_1637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2898;
  reg [31:0] _T_1637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2899;
  reg [31:0] _T_1638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2900;
  reg [31:0] _T_1638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2901;
  reg [31:0] _T_1639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2902;
  reg [31:0] _T_1639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2903;
  reg [31:0] _T_1640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2904;
  reg [31:0] _T_1640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2905;
  reg [31:0] _T_1641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2906;
  reg [31:0] _T_1641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2907;
  reg [31:0] _T_1642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2908;
  reg [31:0] _T_1642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2909;
  reg [31:0] _T_1643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2910;
  reg [31:0] _T_1643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2911;
  reg [31:0] _T_1644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2912;
  reg [31:0] _T_1644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2913;
  reg [31:0] _T_1645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2914;
  reg [31:0] _T_1645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2915;
  reg [31:0] _T_1646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2916;
  reg [31:0] _T_1646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2917;
  reg [31:0] _T_1647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2918;
  reg [31:0] _T_1647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2919;
  reg [31:0] _T_1648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2920;
  reg [31:0] _T_1648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2921;
  reg [31:0] _T_1649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2922;
  reg [31:0] _T_1649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2923;
  reg [31:0] _T_1650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2924;
  reg [31:0] _T_1650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2925;
  reg [31:0] _T_1651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2926;
  reg [31:0] _T_1651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2927;
  reg [31:0] _T_1652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2928;
  reg [31:0] _T_1652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2929;
  reg [31:0] _T_1653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2930;
  reg [31:0] _T_1653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2931;
  reg [31:0] _T_1654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2932;
  reg [31:0] _T_1654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2933;
  reg [31:0] _T_1655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2934;
  reg [31:0] _T_1655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2935;
  reg [31:0] _T_1656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2936;
  reg [31:0] _T_1656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2937;
  reg [31:0] _T_1657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2938;
  reg [31:0] _T_1657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2939;
  reg [31:0] _T_1658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2940;
  reg [31:0] _T_1658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2941;
  reg [31:0] _T_1659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2942;
  reg [31:0] _T_1659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2943;
  reg [31:0] _T_1660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2944;
  reg [31:0] _T_1660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2945;
  reg [31:0] _T_1661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2946;
  reg [31:0] _T_1661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2947;
  reg [31:0] _T_1662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2948;
  reg [31:0] _T_1662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2949;
  reg [31:0] _T_1663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2950;
  reg [31:0] _T_1663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2951;
  reg [31:0] _T_1664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2952;
  reg [31:0] _T_1664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2953;
  reg [31:0] _T_1665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2954;
  reg [31:0] _T_1665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2955;
  reg [31:0] _T_1666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2956;
  reg [31:0] _T_1666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2957;
  reg [31:0] _T_1667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2958;
  reg [31:0] _T_1667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2959;
  reg [31:0] _T_1668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2960;
  reg [31:0] _T_1668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2961;
  reg [31:0] _T_1669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2962;
  reg [31:0] _T_1669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2963;
  reg [31:0] _T_1670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2964;
  reg [31:0] _T_1670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2965;
  reg [31:0] _T_1671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2966;
  reg [31:0] _T_1671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2967;
  reg [31:0] _T_1672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2968;
  reg [31:0] _T_1672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2969;
  reg [31:0] _T_1673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2970;
  reg [31:0] _T_1673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2971;
  reg [31:0] _T_1674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2972;
  reg [31:0] _T_1674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2973;
  reg [31:0] _T_1675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2974;
  reg [31:0] _T_1675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2975;
  reg [31:0] _T_1676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2976;
  reg [31:0] _T_1676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2977;
  reg [31:0] _T_1677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2978;
  reg [31:0] _T_1677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2979;
  reg [31:0] _T_1678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2980;
  reg [31:0] _T_1678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2981;
  reg [31:0] _T_1679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2982;
  reg [31:0] _T_1679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2983;
  reg [31:0] _T_1680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2984;
  reg [31:0] _T_1680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2985;
  reg [31:0] _T_1681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2986;
  reg [31:0] _T_1681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2987;
  reg [31:0] _T_1682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2988;
  reg [31:0] _T_1682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2989;
  reg [31:0] _T_1683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2990;
  reg [31:0] _T_1683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2991;
  reg [31:0] _T_1684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2992;
  reg [31:0] _T_1684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2993;
  reg [31:0] _T_1685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2994;
  reg [31:0] _T_1685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2995;
  reg [31:0] _T_1686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2996;
  reg [31:0] _T_1686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2997;
  reg [31:0] _T_1687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2998;
  reg [31:0] _T_1687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2999;
  reg [31:0] _T_1688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3000;
  reg [31:0] _T_1688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3001;
  reg [31:0] _T_1689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3002;
  reg [31:0] _T_1689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3003;
  reg [31:0] _T_1690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3004;
  reg [31:0] _T_1690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3005;
  reg [31:0] _T_1691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3006;
  reg [31:0] _T_1691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3007;
  reg [31:0] _T_1692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3008;
  reg [31:0] _T_1692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3009;
  reg [31:0] _T_1693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3010;
  reg [31:0] _T_1693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3011;
  reg [31:0] _T_1694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3012;
  reg [31:0] _T_1694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3013;
  reg [31:0] _T_1695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3014;
  reg [31:0] _T_1695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3015;
  reg [31:0] _T_1696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3016;
  reg [31:0] _T_1696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3017;
  reg [31:0] _T_1697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3018;
  reg [31:0] _T_1697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3019;
  reg [31:0] _T_1698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3020;
  reg [31:0] _T_1698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3021;
  reg [31:0] _T_1699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3022;
  reg [31:0] _T_1699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3023;
  reg [31:0] _T_1700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3024;
  reg [31:0] _T_1700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3025;
  reg [31:0] _T_1701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3026;
  reg [31:0] _T_1701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3027;
  reg [31:0] _T_1702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3028;
  reg [31:0] _T_1702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3029;
  reg [31:0] _T_1703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3030;
  reg [31:0] _T_1703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3031;
  reg [31:0] _T_1704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3032;
  reg [31:0] _T_1704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3033;
  reg [31:0] _T_1705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3034;
  reg [31:0] _T_1705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3035;
  reg [31:0] _T_1706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3036;
  reg [31:0] _T_1706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3037;
  reg [31:0] _T_1707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3038;
  reg [31:0] _T_1707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3039;
  reg [31:0] _T_1708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3040;
  reg [31:0] _T_1708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3041;
  reg [31:0] _T_1709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3042;
  reg [31:0] _T_1709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3043;
  reg [31:0] _T_1710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3044;
  reg [31:0] _T_1710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3045;
  reg [31:0] _T_1711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3046;
  reg [31:0] _T_1711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3047;
  reg [31:0] _T_1712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3048;
  reg [31:0] _T_1712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3049;
  reg [31:0] _T_1713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3050;
  reg [31:0] _T_1713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3051;
  reg [31:0] _T_1714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3052;
  reg [31:0] _T_1714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3053;
  reg [31:0] _T_1715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3054;
  reg [31:0] _T_1715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3055;
  reg [31:0] _T_1716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3056;
  reg [31:0] _T_1716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3057;
  reg [31:0] _T_1717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3058;
  reg [31:0] _T_1717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3059;
  reg [31:0] _T_1718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3060;
  reg [31:0] _T_1718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3061;
  reg [31:0] _T_1719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3062;
  reg [31:0] _T_1719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3063;
  reg [31:0] _T_1720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3064;
  reg [31:0] _T_1720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3065;
  reg [31:0] _T_1721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3066;
  reg [31:0] _T_1721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3067;
  reg [31:0] _T_1722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3068;
  reg [31:0] _T_1722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3069;
  reg [31:0] _T_1723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3070;
  reg [31:0] _T_1723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3071;
  reg [31:0] _T_1724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3072;
  reg [31:0] _T_1724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3073;
  reg [31:0] _T_1725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3074;
  reg [31:0] _T_1725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3075;
  reg [31:0] _T_1726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3076;
  reg [31:0] _T_1726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3077;
  reg [31:0] _T_1727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3078;
  reg [31:0] _T_1727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3079;
  reg [31:0] _T_1728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3080;
  reg [31:0] _T_1728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3081;
  reg [31:0] _T_1729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3082;
  reg [31:0] _T_1729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3083;
  reg [31:0] _T_1730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3084;
  reg [31:0] _T_1730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3085;
  reg [31:0] _T_1731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3086;
  reg [31:0] _T_1731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3087;
  reg [31:0] _T_1732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3088;
  reg [31:0] _T_1732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3089;
  reg [31:0] _T_1733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3090;
  reg [31:0] _T_1733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3091;
  reg [31:0] _T_1734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3092;
  reg [31:0] _T_1734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3093;
  reg [31:0] _T_1735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3094;
  reg [31:0] _T_1735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3095;
  reg [31:0] _T_1736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3096;
  reg [31:0] _T_1736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3097;
  reg [31:0] _T_1737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3098;
  reg [31:0] _T_1737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3099;
  reg [31:0] _T_1738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3100;
  reg [31:0] _T_1738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3101;
  reg [31:0] _T_1739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3102;
  reg [31:0] _T_1739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3103;
  reg [31:0] _T_1740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3104;
  reg [31:0] _T_1740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3105;
  reg [31:0] _T_1741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3106;
  reg [31:0] _T_1741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3107;
  reg [31:0] _T_1742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3108;
  reg [31:0] _T_1742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3109;
  reg [31:0] _T_1743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3110;
  reg [31:0] _T_1743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3111;
  reg [31:0] _T_1744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3112;
  reg [31:0] _T_1744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3113;
  reg [31:0] _T_1745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3114;
  reg [31:0] _T_1745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3115;
  reg [31:0] _T_1746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3116;
  reg [31:0] _T_1746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3117;
  reg [31:0] _T_1747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3118;
  reg [31:0] _T_1747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3119;
  reg [31:0] _T_1748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3120;
  reg [31:0] _T_1748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3121;
  reg [31:0] _T_1749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3122;
  reg [31:0] _T_1749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3123;
  reg [31:0] _T_1750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3124;
  reg [31:0] _T_1750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3125;
  reg [31:0] _T_1751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3126;
  reg [31:0] _T_1751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3127;
  reg [31:0] _T_1752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3128;
  reg [31:0] _T_1752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3129;
  reg [31:0] _T_1753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3130;
  reg [31:0] _T_1753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3131;
  reg [31:0] _T_1754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3132;
  reg [31:0] _T_1754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3133;
  reg [31:0] _T_1755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3134;
  reg [31:0] _T_1755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3135;
  reg [31:0] _T_1756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3136;
  reg [31:0] _T_1756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3137;
  reg [31:0] _T_1757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3138;
  reg [31:0] _T_1757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3139;
  reg [31:0] _T_1758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3140;
  reg [31:0] _T_1758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3141;
  reg [31:0] _T_1759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3142;
  reg [31:0] _T_1759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3143;
  reg [31:0] _T_1760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3144;
  reg [31:0] _T_1760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3145;
  reg [31:0] _T_1761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3146;
  reg [31:0] _T_1761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3147;
  reg [31:0] _T_1762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3148;
  reg [31:0] _T_1762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3149;
  reg [31:0] _T_1763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3150;
  reg [31:0] _T_1763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3151;
  reg [31:0] _T_1764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3152;
  reg [31:0] _T_1764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3153;
  reg [31:0] _T_1765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3154;
  reg [31:0] _T_1765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3155;
  reg [31:0] _T_1766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3156;
  reg [31:0] _T_1766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3157;
  reg [31:0] _T_1767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3158;
  reg [31:0] _T_1767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3159;
  reg [31:0] _T_1768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3160;
  reg [31:0] _T_1768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3161;
  reg [31:0] _T_1769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3162;
  reg [31:0] _T_1769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3163;
  reg [31:0] _T_1770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3164;
  reg [31:0] _T_1770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3165;
  reg [31:0] _T_1771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3166;
  reg [31:0] _T_1771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3167;
  reg [31:0] _T_1772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3168;
  reg [31:0] _T_1772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3169;
  reg [31:0] _T_1773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3170;
  reg [31:0] _T_1773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3171;
  reg [31:0] _T_1774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3172;
  reg [31:0] _T_1774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3173;
  reg [31:0] _T_1775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3174;
  reg [31:0] _T_1775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3175;
  reg [31:0] _T_1776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3176;
  reg [31:0] _T_1776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3177;
  reg [31:0] _T_1777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3178;
  reg [31:0] _T_1777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3179;
  reg [31:0] _T_1778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3180;
  reg [31:0] _T_1778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3181;
  reg [31:0] _T_1779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3182;
  reg [31:0] _T_1779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3183;
  reg [31:0] _T_1780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3184;
  reg [31:0] _T_1780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3185;
  reg [31:0] _T_1781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3186;
  reg [31:0] _T_1781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3187;
  reg [31:0] _T_1782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3188;
  reg [31:0] _T_1782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3189;
  reg [31:0] _T_1783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3190;
  reg [31:0] _T_1783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3191;
  reg [31:0] _T_1784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3192;
  reg [31:0] _T_1784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3193;
  reg [31:0] _T_1785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3194;
  reg [31:0] _T_1785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3195;
  reg [31:0] _T_1786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3196;
  reg [31:0] _T_1786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3197;
  reg [31:0] _T_1787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3198;
  reg [31:0] _T_1787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3199;
  reg [31:0] _T_1788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3200;
  reg [31:0] _T_1788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3201;
  reg [31:0] _T_1789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3202;
  reg [31:0] _T_1789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3203;
  reg [31:0] _T_1790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3204;
  reg [31:0] _T_1790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3205;
  reg [31:0] _T_1791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3206;
  reg [31:0] _T_1791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3207;
  reg [31:0] _T_1792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3208;
  reg [31:0] _T_1792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3209;
  reg [31:0] _T_1793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3210;
  reg [31:0] _T_1793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3211;
  reg [31:0] _T_1794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3212;
  reg [31:0] _T_1794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3213;
  reg [31:0] _T_1795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3214;
  reg [31:0] _T_1795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3215;
  reg [31:0] _T_1796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3216;
  reg [31:0] _T_1796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3217;
  reg [31:0] _T_1797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3218;
  reg [31:0] _T_1797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3219;
  reg [31:0] _T_1798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3220;
  reg [31:0] _T_1798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3221;
  reg [31:0] _T_1799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3222;
  reg [31:0] _T_1799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3223;
  reg [31:0] _T_1800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3224;
  reg [31:0] _T_1800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3225;
  reg [31:0] _T_1801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3226;
  reg [31:0] _T_1801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3227;
  reg [31:0] _T_1802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3228;
  reg [31:0] _T_1802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3229;
  reg [31:0] _T_1803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3230;
  reg [31:0] _T_1803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3231;
  reg [31:0] _T_1804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3232;
  reg [31:0] _T_1804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3233;
  reg [31:0] _T_1805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3234;
  reg [31:0] _T_1805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3235;
  reg [31:0] _T_1806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3236;
  reg [31:0] _T_1806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3237;
  reg [31:0] _T_1807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3238;
  reg [31:0] _T_1807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3239;
  reg [31:0] _T_1808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3240;
  reg [31:0] _T_1808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3241;
  reg [31:0] _T_1809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3242;
  reg [31:0] _T_1809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3243;
  reg [31:0] _T_1810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3244;
  reg [31:0] _T_1810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3245;
  reg [31:0] _T_1811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3246;
  reg [31:0] _T_1811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3247;
  reg [31:0] _T_1812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3248;
  reg [31:0] _T_1812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3249;
  reg [31:0] _T_1813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3250;
  reg [31:0] _T_1813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3251;
  reg [31:0] _T_1814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3252;
  reg [31:0] _T_1814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3253;
  reg [31:0] _T_1815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3254;
  reg [31:0] _T_1815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3255;
  reg [31:0] _T_1816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3256;
  reg [31:0] _T_1816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3257;
  reg [31:0] _T_1817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3258;
  reg [31:0] _T_1817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3259;
  reg [31:0] _T_1818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3260;
  reg [31:0] _T_1818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3261;
  reg [31:0] _T_1819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3262;
  reg [31:0] _T_1819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3263;
  reg [31:0] _T_1820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3264;
  reg [31:0] _T_1820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3265;
  reg [31:0] _T_1821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3266;
  reg [31:0] _T_1821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3267;
  reg [31:0] _T_1822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3268;
  reg [31:0] _T_1822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3269;
  reg [31:0] _T_1823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3270;
  reg [31:0] _T_1823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3271;
  reg [31:0] _T_1824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3272;
  reg [31:0] _T_1824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3273;
  reg [31:0] _T_1825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3274;
  reg [31:0] _T_1825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3275;
  reg [31:0] _T_1826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3276;
  reg [31:0] _T_1826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3277;
  reg [31:0] _T_1827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3278;
  reg [31:0] _T_1827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3279;
  reg [31:0] _T_1828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3280;
  reg [31:0] _T_1828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3281;
  reg [31:0] _T_1829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3282;
  reg [31:0] _T_1829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3283;
  reg [31:0] _T_1830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3284;
  reg [31:0] _T_1830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3285;
  reg [31:0] _T_1831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3286;
  reg [31:0] _T_1831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3287;
  reg [31:0] _T_1832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3288;
  reg [31:0] _T_1832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3289;
  reg [31:0] _T_1833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3290;
  reg [31:0] _T_1833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3291;
  reg [31:0] _T_1834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3292;
  reg [31:0] _T_1834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3293;
  reg [31:0] _T_1835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3294;
  reg [31:0] _T_1835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3295;
  reg [31:0] _T_1836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3296;
  reg [31:0] _T_1836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3297;
  reg [31:0] _T_1837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3298;
  reg [31:0] _T_1837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3299;
  reg [31:0] _T_1838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3300;
  reg [31:0] _T_1838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3301;
  reg [31:0] _T_1839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3302;
  reg [31:0] _T_1839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3303;
  reg [31:0] _T_1840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3304;
  reg [31:0] _T_1840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3305;
  reg [31:0] _T_1841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3306;
  reg [31:0] _T_1841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3307;
  reg [31:0] _T_1842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3308;
  reg [31:0] _T_1842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3309;
  reg [31:0] _T_1843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3310;
  reg [31:0] _T_1843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3311;
  reg [31:0] _T_1844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3312;
  reg [31:0] _T_1844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3313;
  reg [31:0] _T_1845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3314;
  reg [31:0] _T_1845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3315;
  reg [31:0] _T_1846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3316;
  reg [31:0] _T_1846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3317;
  reg [31:0] _T_1847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3318;
  reg [31:0] _T_1847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3319;
  reg [31:0] _T_1848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3320;
  reg [31:0] _T_1848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3321;
  reg [31:0] _T_1849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3322;
  reg [31:0] _T_1849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3323;
  reg [31:0] _T_1850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3324;
  reg [31:0] _T_1850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3325;
  reg [31:0] _T_1851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3326;
  reg [31:0] _T_1851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3327;
  reg [31:0] _T_1852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3328;
  reg [31:0] _T_1852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3329;
  reg [31:0] _T_1853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3330;
  reg [31:0] _T_1853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3331;
  reg [31:0] _T_1854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3332;
  reg [31:0] _T_1854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3333;
  reg [31:0] _T_1855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3334;
  reg [31:0] _T_1855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3335;
  reg [31:0] _T_1856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3336;
  reg [31:0] _T_1856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3337;
  reg [31:0] _T_1857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3338;
  reg [31:0] _T_1857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3339;
  reg [31:0] _T_1858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3340;
  reg [31:0] _T_1858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3341;
  reg [31:0] _T_1859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3342;
  reg [31:0] _T_1859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3343;
  reg [31:0] _T_1860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3344;
  reg [31:0] _T_1860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3345;
  reg [31:0] _T_1861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3346;
  reg [31:0] _T_1861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3347;
  reg [31:0] _T_1862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3348;
  reg [31:0] _T_1862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3349;
  reg [31:0] _T_1863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3350;
  reg [31:0] _T_1863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3351;
  reg [31:0] _T_1864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3352;
  reg [31:0] _T_1864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3353;
  reg [31:0] _T_1865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3354;
  reg [31:0] _T_1865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3355;
  reg [31:0] _T_1866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3356;
  reg [31:0] _T_1866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3357;
  reg [31:0] _T_1867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3358;
  reg [31:0] _T_1867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3359;
  reg [31:0] _T_1868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3360;
  reg [31:0] _T_1868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3361;
  reg [31:0] _T_1869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3362;
  reg [31:0] _T_1869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3363;
  reg [31:0] _T_1870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3364;
  reg [31:0] _T_1870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3365;
  reg [31:0] _T_1871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3366;
  reg [31:0] _T_1871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3367;
  reg [31:0] _T_1872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3368;
  reg [31:0] _T_1872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3369;
  reg [31:0] _T_1873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3370;
  reg [31:0] _T_1873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3371;
  reg [31:0] _T_1874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3372;
  reg [31:0] _T_1874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3373;
  reg [31:0] _T_1875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3374;
  reg [31:0] _T_1875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3375;
  reg [31:0] _T_1876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3376;
  reg [31:0] _T_1876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3377;
  reg [31:0] _T_1877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3378;
  reg [31:0] _T_1877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3379;
  reg [31:0] _T_1878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3380;
  reg [31:0] _T_1878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3381;
  reg [31:0] _T_1879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3382;
  reg [31:0] _T_1879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3383;
  reg [31:0] _T_1880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3384;
  reg [31:0] _T_1880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3385;
  reg [31:0] _T_1881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3386;
  reg [31:0] _T_1881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3387;
  reg [31:0] _T_1882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3388;
  reg [31:0] _T_1882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3389;
  reg [31:0] _T_1883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3390;
  reg [31:0] _T_1883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3391;
  reg [31:0] _T_1884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3392;
  reg [31:0] _T_1884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3393;
  reg [31:0] _T_1885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3394;
  reg [31:0] _T_1885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3395;
  reg [31:0] _T_1886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3396;
  reg [31:0] _T_1886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3397;
  reg [31:0] _T_1887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3398;
  reg [31:0] _T_1887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3399;
  reg [31:0] _T_1888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3400;
  reg [31:0] _T_1888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3401;
  reg [31:0] _T_1889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3402;
  reg [31:0] _T_1889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3403;
  reg [31:0] _T_1890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3404;
  reg [31:0] _T_1890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3405;
  reg [31:0] _T_1891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3406;
  reg [31:0] _T_1891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3407;
  reg [31:0] _T_1892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3408;
  reg [31:0] _T_1892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3409;
  reg [31:0] _T_1893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3410;
  reg [31:0] _T_1893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3411;
  reg [31:0] _T_1894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3412;
  reg [31:0] _T_1894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3413;
  reg [31:0] _T_1895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3414;
  reg [31:0] _T_1895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3415;
  reg [31:0] _T_1896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3416;
  reg [31:0] _T_1896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3417;
  reg [31:0] _T_1897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3418;
  reg [31:0] _T_1897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3419;
  reg [31:0] _T_1898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3420;
  reg [31:0] _T_1898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3421;
  reg [31:0] _T_1899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3422;
  reg [31:0] _T_1899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3423;
  reg [31:0] _T_1900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3424;
  reg [31:0] _T_1900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3425;
  reg [31:0] _T_1901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3426;
  reg [31:0] _T_1901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3427;
  reg [31:0] _T_1902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3428;
  reg [31:0] _T_1902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3429;
  reg [31:0] _T_1903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3430;
  reg [31:0] _T_1903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3431;
  reg [31:0] _T_1904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3432;
  reg [31:0] _T_1904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3433;
  reg [31:0] _T_1905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3434;
  reg [31:0] _T_1905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3435;
  reg [31:0] _T_1906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3436;
  reg [31:0] _T_1906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3437;
  reg [31:0] _T_1907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3438;
  reg [31:0] _T_1907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3439;
  reg [31:0] _T_1908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3440;
  reg [31:0] _T_1908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3441;
  reg [31:0] _T_1909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3442;
  reg [31:0] _T_1909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3443;
  reg [31:0] _T_1910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3444;
  reg [31:0] _T_1910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3445;
  reg [31:0] _T_1911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3446;
  reg [31:0] _T_1911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3447;
  reg [31:0] _T_1912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3448;
  reg [31:0] _T_1912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3449;
  reg [31:0] _T_1913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3450;
  reg [31:0] _T_1913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3451;
  reg [31:0] _T_1914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3452;
  reg [31:0] _T_1914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3453;
  reg [31:0] _T_1915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3454;
  reg [31:0] _T_1915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3455;
  reg [31:0] _T_1916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3456;
  reg [31:0] _T_1916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3457;
  reg [31:0] _T_1917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3458;
  reg [31:0] _T_1917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3459;
  reg [31:0] _T_1918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3460;
  reg [31:0] _T_1918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3461;
  reg [31:0] _T_1919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3462;
  reg [31:0] _T_1919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3463;
  reg [31:0] _T_1920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3464;
  reg [31:0] _T_1920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3465;
  reg [31:0] _T_1921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3466;
  reg [31:0] _T_1921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3467;
  reg [31:0] _T_1922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3468;
  reg [31:0] _T_1922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3469;
  reg [31:0] _T_1923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3470;
  reg [31:0] _T_1923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3471;
  reg [31:0] _T_1924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3472;
  reg [31:0] _T_1924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3473;
  reg [31:0] _T_1925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3474;
  reg [31:0] _T_1925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3475;
  reg [31:0] _T_1926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3476;
  reg [31:0] _T_1926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3477;
  reg [31:0] _T_1927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3478;
  reg [31:0] _T_1927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3479;
  reg [31:0] _T_1928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3480;
  reg [31:0] _T_1928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3481;
  reg [31:0] _T_1929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3482;
  reg [31:0] _T_1929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3483;
  reg [31:0] _T_1930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3484;
  reg [31:0] _T_1930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3485;
  reg [31:0] _T_1931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3486;
  reg [31:0] _T_1931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3487;
  reg [31:0] _T_1932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3488;
  reg [31:0] _T_1932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3489;
  reg [31:0] _T_1933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3490;
  reg [31:0] _T_1933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3491;
  reg [31:0] _T_1934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3492;
  reg [31:0] _T_1934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3493;
  reg [31:0] _T_1935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3494;
  reg [31:0] _T_1935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3495;
  reg [31:0] _T_1936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3496;
  reg [31:0] _T_1936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3497;
  reg [31:0] _T_1937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3498;
  reg [31:0] _T_1937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3499;
  reg [31:0] _T_1938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3500;
  reg [31:0] _T_1938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3501;
  reg [31:0] _T_1939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3502;
  reg [31:0] _T_1939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3503;
  reg [31:0] _T_1940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3504;
  reg [31:0] _T_1940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3505;
  reg [31:0] _T_1941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3506;
  reg [31:0] _T_1941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3507;
  reg [31:0] _T_1942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3508;
  reg [31:0] _T_1942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3509;
  reg [31:0] _T_1943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3510;
  reg [31:0] _T_1943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3511;
  reg [31:0] _T_1944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3512;
  reg [31:0] _T_1944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3513;
  reg [31:0] _T_1945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3514;
  reg [31:0] _T_1945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3515;
  reg [31:0] _T_1946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3516;
  reg [31:0] _T_1946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3517;
  reg [31:0] _T_1947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3518;
  reg [31:0] _T_1947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3519;
  reg [31:0] _T_1948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3520;
  reg [31:0] _T_1948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3521;
  reg [31:0] _T_1949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3522;
  reg [31:0] _T_1949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3523;
  reg [31:0] _T_1950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3524;
  reg [31:0] _T_1950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3525;
  reg [31:0] _T_1951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3526;
  reg [31:0] _T_1951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3527;
  reg [31:0] _T_1952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3528;
  reg [31:0] _T_1952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3529;
  reg [31:0] _T_1953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3530;
  reg [31:0] _T_1953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3531;
  reg [31:0] _T_1954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3532;
  reg [31:0] _T_1954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3533;
  reg [31:0] _T_1955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3534;
  reg [31:0] _T_1955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3535;
  reg [31:0] _T_1956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3536;
  reg [31:0] _T_1956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3537;
  reg [31:0] _T_1957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3538;
  reg [31:0] _T_1957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3539;
  reg [31:0] _T_1958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3540;
  reg [31:0] _T_1958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3541;
  reg [31:0] _T_1959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3542;
  reg [31:0] _T_1959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3543;
  reg [31:0] _T_1960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3544;
  reg [31:0] _T_1960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3545;
  reg [31:0] _T_1961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3546;
  reg [31:0] _T_1961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3547;
  reg [31:0] _T_1962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3548;
  reg [31:0] _T_1962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3549;
  reg [31:0] _T_1963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3550;
  reg [31:0] _T_1963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3551;
  reg [31:0] _T_1964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3552;
  reg [31:0] _T_1964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3553;
  reg [31:0] _T_1965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3554;
  reg [31:0] _T_1965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3555;
  reg [31:0] _T_1966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3556;
  reg [31:0] _T_1966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3557;
  reg [31:0] _T_1967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3558;
  reg [31:0] _T_1967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3559;
  reg [31:0] _T_1968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3560;
  reg [31:0] _T_1968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3561;
  reg [31:0] _T_1969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3562;
  reg [31:0] _T_1969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3563;
  reg [31:0] _T_1970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3564;
  reg [31:0] _T_1970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3565;
  reg [31:0] _T_1971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3566;
  reg [31:0] _T_1971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3567;
  reg [31:0] _T_1972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3568;
  reg [31:0] _T_1972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3569;
  reg [31:0] _T_1973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3570;
  reg [31:0] _T_1973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3571;
  reg [31:0] _T_1974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3572;
  reg [31:0] _T_1974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3573;
  reg [31:0] _T_1975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3574;
  reg [31:0] _T_1975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3575;
  reg [31:0] _T_1976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3576;
  reg [31:0] _T_1976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3577;
  reg [31:0] _T_1977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3578;
  reg [31:0] _T_1977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3579;
  reg [31:0] _T_1978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3580;
  reg [31:0] _T_1978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3581;
  reg [31:0] _T_1979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3582;
  reg [31:0] _T_1979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3583;
  reg [31:0] _T_1980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3584;
  reg [31:0] _T_1980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3585;
  reg [31:0] _T_1981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3586;
  reg [31:0] _T_1981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3587;
  reg [31:0] _T_1982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3588;
  reg [31:0] _T_1982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3589;
  reg [31:0] _T_1983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3590;
  reg [31:0] _T_1983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3591;
  reg [31:0] _T_1984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3592;
  reg [31:0] _T_1984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3593;
  reg [31:0] _T_1985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3594;
  reg [31:0] _T_1985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3595;
  reg [31:0] _T_1986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3596;
  reg [31:0] _T_1986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3597;
  reg [31:0] _T_1987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3598;
  reg [31:0] _T_1987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3599;
  reg [31:0] _T_1988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3600;
  reg [31:0] _T_1988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3601;
  reg [31:0] _T_1989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3602;
  reg [31:0] _T_1989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3603;
  reg [31:0] _T_1990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3604;
  reg [31:0] _T_1990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3605;
  reg [31:0] _T_1991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3606;
  reg [31:0] _T_1991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3607;
  reg [31:0] _T_1992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3608;
  reg [31:0] _T_1992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3609;
  reg [31:0] _T_1993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3610;
  reg [31:0] _T_1993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3611;
  reg [31:0] _T_1994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3612;
  reg [31:0] _T_1994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3613;
  reg [31:0] _T_1995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3614;
  reg [31:0] _T_1995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3615;
  reg [31:0] _T_1996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3616;
  reg [31:0] _T_1996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3617;
  reg [31:0] _T_1997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3618;
  reg [31:0] _T_1997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3619;
  reg [31:0] _T_1998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3620;
  reg [31:0] _T_1998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3621;
  reg [31:0] _T_1999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3622;
  reg [31:0] _T_1999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3623;
  reg [31:0] _T_2000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3624;
  reg [31:0] _T_2000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3625;
  reg [31:0] _T_2001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3626;
  reg [31:0] _T_2001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3627;
  reg [31:0] _T_2002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3628;
  reg [31:0] _T_2002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3629;
  reg [31:0] _T_2003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3630;
  reg [31:0] _T_2003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3631;
  reg [31:0] _T_2004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3632;
  reg [31:0] _T_2004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3633;
  reg [31:0] _T_2005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3634;
  reg [31:0] _T_2005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3635;
  reg [31:0] _T_2006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3636;
  reg [31:0] _T_2006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3637;
  reg [31:0] _T_2007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3638;
  reg [31:0] _T_2007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3639;
  reg [31:0] _T_2008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3640;
  reg [31:0] _T_2008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3641;
  reg [31:0] _T_2009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3642;
  reg [31:0] _T_2009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3643;
  reg [31:0] _T_2010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3644;
  reg [31:0] _T_2010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3645;
  reg [31:0] _T_2011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3646;
  reg [31:0] _T_2011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3647;
  reg [31:0] _T_2012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3648;
  reg [31:0] _T_2012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3649;
  reg [31:0] _T_2013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3650;
  reg [31:0] _T_2013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3651;
  reg [31:0] _T_2014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3652;
  reg [31:0] _T_2014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3653;
  reg [31:0] _T_2015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3654;
  reg [31:0] _T_2015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3655;
  reg [31:0] _T_2016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3656;
  reg [31:0] _T_2016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3657;
  reg [31:0] _T_2017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3658;
  reg [31:0] _T_2017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3659;
  reg [31:0] _T_2018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3660;
  reg [31:0] _T_2018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3661;
  reg [31:0] _T_2019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3662;
  reg [31:0] _T_2019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3663;
  reg [31:0] _T_2020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3664;
  reg [31:0] _T_2020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3665;
  reg [31:0] _T_2021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3666;
  reg [31:0] _T_2021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3667;
  reg [31:0] _T_2022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3668;
  reg [31:0] _T_2022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3669;
  reg [31:0] _T_2023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3670;
  reg [31:0] _T_2023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3671;
  reg [31:0] _T_2024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3672;
  reg [31:0] _T_2024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3673;
  reg [31:0] _T_2025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3674;
  reg [31:0] _T_2025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3675;
  reg [31:0] _T_2026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3676;
  reg [31:0] _T_2026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3677;
  reg [31:0] _T_2027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3678;
  reg [31:0] _T_2027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3679;
  reg [31:0] _T_2028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3680;
  reg [31:0] _T_2028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3681;
  reg [31:0] _T_2029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3682;
  reg [31:0] _T_2029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3683;
  reg [31:0] _T_2030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3684;
  reg [31:0] _T_2030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3685;
  reg [31:0] _T_2031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3686;
  reg [31:0] _T_2031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3687;
  reg [31:0] _T_2032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3688;
  reg [31:0] _T_2032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3689;
  reg [31:0] _T_2033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3690;
  reg [31:0] _T_2033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3691;
  reg [31:0] _T_2034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3692;
  reg [31:0] _T_2034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3693;
  reg [31:0] _T_2035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3694;
  reg [31:0] _T_2035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3695;
  reg [31:0] _T_2036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3696;
  reg [31:0] _T_2036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3697;
  reg [31:0] _T_2037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3698;
  reg [31:0] _T_2037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3699;
  reg [31:0] _T_2038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3700;
  reg [31:0] _T_2038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3701;
  reg [31:0] _T_2039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3702;
  reg [31:0] _T_2039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3703;
  reg [31:0] _T_2040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3704;
  reg [31:0] _T_2040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3705;
  reg [31:0] _T_2041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3706;
  reg [31:0] _T_2041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3707;
  reg [31:0] _T_2042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3708;
  reg [31:0] _T_2042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3709;
  reg [31:0] _T_2043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3710;
  reg [31:0] _T_2043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3711;
  reg [31:0] _T_2044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3712;
  reg [31:0] _T_2044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3713;
  reg [31:0] _T_2045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3714;
  reg [31:0] _T_2045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3715;
  reg [31:0] _T_2046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3716;
  reg [31:0] _T_2046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3717;
  reg [31:0] _T_2047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3718;
  reg [31:0] _T_2047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3719;
  reg [31:0] _T_2048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3720;
  reg [31:0] _T_2048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3721;
  reg [31:0] _T_2049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3722;
  reg [31:0] _T_2049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3723;
  reg [31:0] _T_2050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3724;
  reg [31:0] _T_2050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3725;
  reg [31:0] _T_2051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3726;
  reg [31:0] _T_2051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3727;
  reg [31:0] _T_2052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3728;
  reg [31:0] _T_2052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3729;
  reg [31:0] _T_2053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3730;
  reg [31:0] _T_2053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3731;
  reg [31:0] _T_2054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3732;
  reg [31:0] _T_2054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3733;
  reg [31:0] _T_2055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3734;
  reg [31:0] _T_2055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3735;
  reg [31:0] _T_2056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3736;
  reg [31:0] _T_2056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3737;
  reg [31:0] _T_2057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3738;
  reg [31:0] _T_2057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3739;
  reg [31:0] _T_2058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3740;
  reg [31:0] _T_2058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3741;
  reg [31:0] _T_2059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3742;
  reg [31:0] _T_2059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3743;
  reg [31:0] _T_2060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3744;
  reg [31:0] _T_2060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3745;
  reg [31:0] _T_2061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3746;
  reg [31:0] _T_2061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3747;
  reg [31:0] _T_2062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3748;
  reg [31:0] _T_2062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3749;
  reg [31:0] _T_2063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3750;
  reg [31:0] _T_2063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3751;
  reg [31:0] _T_2064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3752;
  reg [31:0] _T_2064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3753;
  reg [31:0] _T_2065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3754;
  reg [31:0] _T_2065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3755;
  reg [31:0] _T_2066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3756;
  reg [31:0] _T_2066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3757;
  reg [31:0] _T_2067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3758;
  reg [31:0] _T_2067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3759;
  reg [31:0] _T_2068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3760;
  reg [31:0] _T_2068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3761;
  reg [31:0] _T_2069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3762;
  reg [31:0] _T_2069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3763;
  reg [31:0] _T_2070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3764;
  reg [31:0] _T_2070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3765;
  reg [31:0] _T_2071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3766;
  reg [31:0] _T_2071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3767;
  reg [31:0] _T_2072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3768;
  reg [31:0] _T_2072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3769;
  reg [31:0] _T_2073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3770;
  reg [31:0] _T_2073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3771;
  reg [31:0] _T_2074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3772;
  reg [31:0] _T_2074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3773;
  reg [31:0] _T_2075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3774;
  reg [31:0] _T_2075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3775;
  reg [31:0] _T_2076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3776;
  reg [31:0] _T_2076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3777;
  reg [31:0] _T_2077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3778;
  reg [31:0] _T_2077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3779;
  reg [31:0] _T_2078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3780;
  reg [31:0] _T_2078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3781;
  reg [31:0] _T_2079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3782;
  reg [31:0] _T_2079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3783;
  reg [31:0] _T_2080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3784;
  reg [31:0] _T_2080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3785;
  reg [31:0] _T_2081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3786;
  reg [31:0] _T_2081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3787;
  reg [31:0] _T_2082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3788;
  reg [31:0] _T_2082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3789;
  reg [31:0] _T_2083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3790;
  reg [31:0] _T_2083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3791;
  reg [31:0] _T_2084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3792;
  reg [31:0] _T_2084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3793;
  reg [31:0] _T_2085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3794;
  reg [31:0] _T_2085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3795;
  reg [31:0] _T_2086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3796;
  reg [31:0] _T_2086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3797;
  reg [31:0] _T_2087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3798;
  reg [31:0] _T_2087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3799;
  reg [31:0] _T_2088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3800;
  reg [31:0] _T_2088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3801;
  reg [31:0] _T_2089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3802;
  reg [31:0] _T_2089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3803;
  reg [31:0] _T_2090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3804;
  reg [31:0] _T_2090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3805;
  reg [31:0] _T_2091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3806;
  reg [31:0] _T_2091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3807;
  reg [31:0] _T_2092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3808;
  reg [31:0] _T_2092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3809;
  reg [31:0] _T_2093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3810;
  reg [31:0] _T_2093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3811;
  reg [31:0] _T_2094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3812;
  reg [31:0] _T_2094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3813;
  reg [31:0] _T_2095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3814;
  reg [31:0] _T_2095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3815;
  reg [31:0] _T_2096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3816;
  reg [31:0] _T_2096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3817;
  reg [31:0] _T_2097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3818;
  reg [31:0] _T_2097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3819;
  reg [31:0] _T_2098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3820;
  reg [31:0] _T_2098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3821;
  reg [31:0] _T_2099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3822;
  reg [31:0] _T_2099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3823;
  reg [31:0] _T_2100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3824;
  reg [31:0] _T_2100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3825;
  reg [31:0] _T_2101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3826;
  reg [31:0] _T_2101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3827;
  reg [31:0] _T_2102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3828;
  reg [31:0] _T_2102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3829;
  reg [31:0] _T_2103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3830;
  reg [31:0] _T_2103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3831;
  reg [31:0] _T_2104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3832;
  reg [31:0] _T_2104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3833;
  reg [31:0] _T_2105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3834;
  reg [31:0] _T_2105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3835;
  reg [31:0] _T_2106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3836;
  reg [31:0] _T_2106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3837;
  reg [31:0] _T_2107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3838;
  reg [31:0] _T_2107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3839;
  reg [31:0] _T_2108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3840;
  reg [31:0] _T_2108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3841;
  reg [31:0] _T_2109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3842;
  reg [31:0] _T_2109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3843;
  reg [31:0] _T_2110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3844;
  reg [31:0] _T_2110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3845;
  reg [31:0] _T_2111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3846;
  reg [31:0] _T_2111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3847;
  reg [31:0] _T_2112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3848;
  reg [31:0] _T_2112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3849;
  reg [31:0] _T_2113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3850;
  reg [31:0] _T_2113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3851;
  reg [31:0] _T_2114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3852;
  reg [31:0] _T_2114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3853;
  reg [31:0] _T_2115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3854;
  reg [31:0] _T_2115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3855;
  reg [31:0] _T_2116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3856;
  reg [31:0] _T_2116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3857;
  reg [31:0] _T_2117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3858;
  reg [31:0] _T_2117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3859;
  reg [31:0] _T_2118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3860;
  reg [31:0] _T_2118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3861;
  reg [31:0] _T_2119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3862;
  reg [31:0] _T_2119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3863;
  reg [31:0] _T_2120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3864;
  reg [31:0] _T_2120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3865;
  reg [31:0] _T_2121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3866;
  reg [31:0] _T_2121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3867;
  reg [31:0] _T_2122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3868;
  reg [31:0] _T_2122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3869;
  reg [31:0] _T_2123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3870;
  reg [31:0] _T_2123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3871;
  reg [31:0] _T_2124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3872;
  reg [31:0] _T_2124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3873;
  reg [31:0] _T_2125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3874;
  reg [31:0] _T_2125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3875;
  reg [31:0] _T_2126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3876;
  reg [31:0] _T_2126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3877;
  reg [31:0] _T_2127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3878;
  reg [31:0] _T_2127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3879;
  reg [31:0] _T_2128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3880;
  reg [31:0] _T_2128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3881;
  reg [31:0] _T_2129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3882;
  reg [31:0] _T_2129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3883;
  reg [31:0] _T_2130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3884;
  reg [31:0] _T_2130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3885;
  reg [31:0] _T_2131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3886;
  reg [31:0] _T_2131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3887;
  reg [31:0] _T_2132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3888;
  reg [31:0] _T_2132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3889;
  reg [31:0] _T_2133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3890;
  reg [31:0] _T_2133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3891;
  reg [31:0] _T_2134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3892;
  reg [31:0] _T_2134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3893;
  reg [31:0] _T_2135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3894;
  reg [31:0] _T_2135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3895;
  reg [31:0] _T_2136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3896;
  reg [31:0] _T_2136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3897;
  reg [31:0] _T_2137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3898;
  reg [31:0] _T_2137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3899;
  reg [31:0] _T_2138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3900;
  reg [31:0] _T_2138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3901;
  reg [31:0] _T_2139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3902;
  reg [31:0] _T_2139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3903;
  reg [31:0] _T_2140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3904;
  reg [31:0] _T_2140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3905;
  reg [31:0] _T_2141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3906;
  reg [31:0] _T_2141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3907;
  reg [31:0] _T_2142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3908;
  reg [31:0] _T_2142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3909;
  reg [31:0] _T_2143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3910;
  reg [31:0] _T_2143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3911;
  reg [31:0] _T_2144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3912;
  reg [31:0] _T_2144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3913;
  reg [31:0] _T_2145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3914;
  reg [31:0] _T_2145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3915;
  reg [31:0] _T_2146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3916;
  reg [31:0] _T_2146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3917;
  reg [31:0] _T_2147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3918;
  reg [31:0] _T_2147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3919;
  reg [31:0] _T_2148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3920;
  reg [31:0] _T_2148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3921;
  reg [31:0] _T_2149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3922;
  reg [31:0] _T_2149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3923;
  reg [31:0] _T_2150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3924;
  reg [31:0] _T_2150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3925;
  reg [31:0] _T_2151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3926;
  reg [31:0] _T_2151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3927;
  reg [31:0] _T_2152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3928;
  reg [31:0] _T_2152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3929;
  reg [31:0] _T_2153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3930;
  reg [31:0] _T_2153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3931;
  reg [31:0] _T_2154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3932;
  reg [31:0] _T_2154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3933;
  reg [31:0] _T_2155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3934;
  reg [31:0] _T_2155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3935;
  reg [31:0] _T_2156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3936;
  reg [31:0] _T_2156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3937;
  reg [31:0] _T_2157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3938;
  reg [31:0] _T_2157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3939;
  reg [31:0] _T_2158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3940;
  reg [31:0] _T_2158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3941;
  reg [31:0] _T_2159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3942;
  reg [31:0] _T_2159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3943;
  reg [31:0] _T_2160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3944;
  reg [31:0] _T_2160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3945;
  reg [31:0] _T_2161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3946;
  reg [31:0] _T_2161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3947;
  reg [31:0] _T_2162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3948;
  reg [31:0] _T_2162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3949;
  reg [31:0] _T_2163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3950;
  reg [31:0] _T_2163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3951;
  reg [31:0] _T_2164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3952;
  reg [31:0] _T_2164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3953;
  reg [31:0] _T_2165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3954;
  reg [31:0] _T_2165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3955;
  reg [31:0] _T_2166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3956;
  reg [31:0] _T_2166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3957;
  reg [31:0] _T_2167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3958;
  reg [31:0] _T_2167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3959;
  reg [31:0] _T_2168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3960;
  reg [31:0] _T_2168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3961;
  reg [31:0] _T_2169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3962;
  reg [31:0] _T_2169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3963;
  reg [31:0] _T_2170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3964;
  reg [31:0] _T_2170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3965;
  reg [31:0] _T_2171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3966;
  reg [31:0] _T_2171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3967;
  reg [31:0] _T_2172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3968;
  reg [31:0] _T_2172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3969;
  reg [31:0] _T_2173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3970;
  reg [31:0] _T_2173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3971;
  reg [31:0] _T_2174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3972;
  reg [31:0] _T_2174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3973;
  reg [31:0] _T_2175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3974;
  reg [31:0] _T_2175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3975;
  reg [31:0] _T_2176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3976;
  reg [31:0] _T_2176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3977;
  reg [31:0] _T_2177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3978;
  reg [31:0] _T_2177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3979;
  reg [31:0] _T_2178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3980;
  reg [31:0] _T_2178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3981;
  reg [31:0] _T_2179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3982;
  reg [31:0] _T_2179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3983;
  reg [31:0] _T_2180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3984;
  reg [31:0] _T_2180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3985;
  reg [31:0] _T_2181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3986;
  reg [31:0] _T_2181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3987;
  reg [31:0] _T_2182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3988;
  reg [31:0] _T_2182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3989;
  reg [31:0] _T_2183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3990;
  reg [31:0] _T_2183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3991;
  reg [31:0] _T_2184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3992;
  reg [31:0] _T_2184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3993;
  reg [31:0] _T_2185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3994;
  reg [31:0] _T_2185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3995;
  reg [31:0] _T_2186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3996;
  reg [31:0] _T_2186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3997;
  reg [31:0] _T_2187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3998;
  reg [31:0] _T_2187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3999;
  reg [31:0] _T_2188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4000;
  reg [31:0] _T_2188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4001;
  reg [31:0] _T_2189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4002;
  reg [31:0] _T_2189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4003;
  reg [31:0] _T_2190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4004;
  reg [31:0] _T_2190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4005;
  reg [31:0] _T_2191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4006;
  reg [31:0] _T_2191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4007;
  reg [31:0] _T_2192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4008;
  reg [31:0] _T_2192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4009;
  reg [31:0] _T_2193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4010;
  reg [31:0] _T_2193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4011;
  reg [31:0] _T_2194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4012;
  reg [31:0] _T_2194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4013;
  reg [31:0] _T_2195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4014;
  reg [31:0] _T_2195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4015;
  reg [31:0] _T_2196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4016;
  reg [31:0] _T_2196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4017;
  reg [31:0] _T_2197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4018;
  reg [31:0] _T_2197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4019;
  reg [31:0] _T_2198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4020;
  reg [31:0] _T_2198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4021;
  reg [31:0] _T_2199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4022;
  reg [31:0] _T_2199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4023;
  reg [31:0] _T_2200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4024;
  reg [31:0] _T_2200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4025;
  reg [31:0] _T_2201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4026;
  reg [31:0] _T_2201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4027;
  reg [31:0] _T_2202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4028;
  reg [31:0] _T_2202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4029;
  reg [31:0] _T_2203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4030;
  reg [31:0] _T_2203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4031;
  reg [31:0] _T_2204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4032;
  reg [31:0] _T_2204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4033;
  reg [31:0] _T_2205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4034;
  reg [31:0] _T_2205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4035;
  reg [31:0] _T_2206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4036;
  reg [31:0] _T_2206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4037;
  reg [31:0] _T_2207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4038;
  reg [31:0] _T_2207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4039;
  reg [31:0] _T_2208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4040;
  reg [31:0] _T_2208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4041;
  reg [31:0] _T_2209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4042;
  reg [31:0] _T_2209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4043;
  reg [31:0] _T_2210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4044;
  reg [31:0] _T_2210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4045;
  reg [31:0] _T_2211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4046;
  reg [31:0] _T_2211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4047;
  reg [31:0] _T_2212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4048;
  reg [31:0] _T_2212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4049;
  reg [31:0] _T_2213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4050;
  reg [31:0] _T_2213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4051;
  reg [31:0] _T_2214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4052;
  reg [31:0] _T_2214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4053;
  reg [31:0] _T_2215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4054;
  reg [31:0] _T_2215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4055;
  reg [31:0] _T_2216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4056;
  reg [31:0] _T_2216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4057;
  reg [31:0] _T_2217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4058;
  reg [31:0] _T_2217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4059;
  reg [31:0] _T_2218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4060;
  reg [31:0] _T_2218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4061;
  reg [31:0] _T_2219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4062;
  reg [31:0] _T_2219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4063;
  reg [31:0] _T_2220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4064;
  reg [31:0] _T_2220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4065;
  reg [31:0] _T_2221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4066;
  reg [31:0] _T_2221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4067;
  reg [31:0] _T_2222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4068;
  reg [31:0] _T_2222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4069;
  reg [31:0] _T_2223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4070;
  reg [31:0] _T_2223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4071;
  reg [31:0] _T_2224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4072;
  reg [31:0] _T_2224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4073;
  reg [31:0] _T_2225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4074;
  reg [31:0] _T_2225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4075;
  reg [31:0] _T_2226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4076;
  reg [31:0] _T_2226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4077;
  reg [31:0] _T_2227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4078;
  reg [31:0] _T_2227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4079;
  reg [31:0] _T_2228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4080;
  reg [31:0] _T_2228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4081;
  reg [31:0] _T_2229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4082;
  reg [31:0] _T_2229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4083;
  reg [31:0] _T_2230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4084;
  reg [31:0] _T_2230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4085;
  reg [31:0] _T_2231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4086;
  reg [31:0] _T_2231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4087;
  reg [31:0] _T_2232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4088;
  reg [31:0] _T_2232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4089;
  reg [31:0] _T_2233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4090;
  reg [31:0] _T_2233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4091;
  reg [31:0] _T_2234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4092;
  reg [31:0] _T_2234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4093;
  reg [31:0] _T_2235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4094;
  reg [31:0] _T_2235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4095;
  reg [31:0] _T_2236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4096;
  reg [31:0] _T_2236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4097;
  reg [31:0] _T_2239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4098;
  reg [31:0] _T_2239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4099;
  reg [31:0] _T_2240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4100;
  reg [31:0] _T_2240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4101;
  reg [31:0] _T_2241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4102;
  reg [31:0] _T_2241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4103;
  reg [31:0] _T_2242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4104;
  reg [31:0] _T_2242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4105;
  reg [31:0] _T_2243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4106;
  reg [31:0] _T_2243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4107;
  reg [31:0] _T_2244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4108;
  reg [31:0] _T_2244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4109;
  reg [31:0] _T_2245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4110;
  reg [31:0] _T_2245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4111;
  reg [31:0] _T_2246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4112;
  reg [31:0] _T_2246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4113;
  reg [31:0] _T_2247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4114;
  reg [31:0] _T_2247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4115;
  reg [31:0] _T_2248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4116;
  reg [31:0] _T_2248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4117;
  reg [31:0] _T_2249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4118;
  reg [31:0] _T_2249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4119;
  reg [31:0] _T_2250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4120;
  reg [31:0] _T_2250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4121;
  reg [31:0] _T_2251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4122;
  reg [31:0] _T_2251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4123;
  reg [31:0] _T_2252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4124;
  reg [31:0] _T_2252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4125;
  reg [31:0] _T_2253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4126;
  reg [31:0] _T_2253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4127;
  reg [31:0] _T_2254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4128;
  reg [31:0] _T_2254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4129;
  reg [31:0] _T_2255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4130;
  reg [31:0] _T_2255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4131;
  reg [31:0] _T_2256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4132;
  reg [31:0] _T_2256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4133;
  reg [31:0] _T_2257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4134;
  reg [31:0] _T_2257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4135;
  reg [31:0] _T_2258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4136;
  reg [31:0] _T_2258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4137;
  reg [31:0] _T_2259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4138;
  reg [31:0] _T_2259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4139;
  reg [31:0] _T_2260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4140;
  reg [31:0] _T_2260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4141;
  reg [31:0] _T_2261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4142;
  reg [31:0] _T_2261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4143;
  reg [31:0] _T_2262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4144;
  reg [31:0] _T_2262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4145;
  reg [31:0] _T_2263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4146;
  reg [31:0] _T_2263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4147;
  reg [31:0] _T_2264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4148;
  reg [31:0] _T_2264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4149;
  reg [31:0] _T_2265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4150;
  reg [31:0] _T_2265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4151;
  reg [31:0] _T_2266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4152;
  reg [31:0] _T_2266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4153;
  reg [31:0] _T_2267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4154;
  reg [31:0] _T_2267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4155;
  reg [31:0] _T_2268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4156;
  reg [31:0] _T_2268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4157;
  reg [31:0] _T_2269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4158;
  reg [31:0] _T_2269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4159;
  reg [31:0] _T_2270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4160;
  reg [31:0] _T_2270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4161;
  reg [31:0] _T_2271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4162;
  reg [31:0] _T_2271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4163;
  reg [31:0] _T_2272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4164;
  reg [31:0] _T_2272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4165;
  reg [31:0] _T_2273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4166;
  reg [31:0] _T_2273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4167;
  reg [31:0] _T_2274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4168;
  reg [31:0] _T_2274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4169;
  reg [31:0] _T_2275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4170;
  reg [31:0] _T_2275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4171;
  reg [31:0] _T_2276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4172;
  reg [31:0] _T_2276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4173;
  reg [31:0] _T_2277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4174;
  reg [31:0] _T_2277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4175;
  reg [31:0] _T_2278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4176;
  reg [31:0] _T_2278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4177;
  reg [31:0] _T_2279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4178;
  reg [31:0] _T_2279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4179;
  reg [31:0] _T_2280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4180;
  reg [31:0] _T_2280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4181;
  reg [31:0] _T_2281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4182;
  reg [31:0] _T_2281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4183;
  reg [31:0] _T_2282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4184;
  reg [31:0] _T_2282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4185;
  reg [31:0] _T_2283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4186;
  reg [31:0] _T_2283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4187;
  reg [31:0] _T_2284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4188;
  reg [31:0] _T_2284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4189;
  reg [31:0] _T_2285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4190;
  reg [31:0] _T_2285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4191;
  reg [31:0] _T_2286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4192;
  reg [31:0] _T_2286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4193;
  reg [31:0] _T_2287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4194;
  reg [31:0] _T_2287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4195;
  reg [31:0] _T_2288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4196;
  reg [31:0] _T_2288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4197;
  reg [31:0] _T_2289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4198;
  reg [31:0] _T_2289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4199;
  reg [31:0] _T_2290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4200;
  reg [31:0] _T_2290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4201;
  reg [31:0] _T_2291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4202;
  reg [31:0] _T_2291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4203;
  reg [31:0] _T_2292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4204;
  reg [31:0] _T_2292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4205;
  reg [31:0] _T_2293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4206;
  reg [31:0] _T_2293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4207;
  reg [31:0] _T_2294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4208;
  reg [31:0] _T_2294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4209;
  reg [31:0] _T_2295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4210;
  reg [31:0] _T_2295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4211;
  reg [31:0] _T_2296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4212;
  reg [31:0] _T_2296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4213;
  reg [31:0] _T_2297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4214;
  reg [31:0] _T_2297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4215;
  reg [31:0] _T_2298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4216;
  reg [31:0] _T_2298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4217;
  reg [31:0] _T_2299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4218;
  reg [31:0] _T_2299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4219;
  reg [31:0] _T_2300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4220;
  reg [31:0] _T_2300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4221;
  reg [31:0] _T_2301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4222;
  reg [31:0] _T_2301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4223;
  reg [31:0] _T_2302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4224;
  reg [31:0] _T_2302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4225;
  reg [31:0] _T_2303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4226;
  reg [31:0] _T_2303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4227;
  reg [31:0] _T_2304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4228;
  reg [31:0] _T_2304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4229;
  reg [31:0] _T_2305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4230;
  reg [31:0] _T_2305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4231;
  reg [31:0] _T_2306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4232;
  reg [31:0] _T_2306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4233;
  reg [31:0] _T_2307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4234;
  reg [31:0] _T_2307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4235;
  reg [31:0] _T_2308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4236;
  reg [31:0] _T_2308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4237;
  reg [31:0] _T_2309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4238;
  reg [31:0] _T_2309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4239;
  reg [31:0] _T_2310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4240;
  reg [31:0] _T_2310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4241;
  reg [31:0] _T_2311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4242;
  reg [31:0] _T_2311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4243;
  reg [31:0] _T_2312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4244;
  reg [31:0] _T_2312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4245;
  reg [31:0] _T_2313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4246;
  reg [31:0] _T_2313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4247;
  reg [31:0] _T_2314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4248;
  reg [31:0] _T_2314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4249;
  reg [31:0] _T_2315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4250;
  reg [31:0] _T_2315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4251;
  reg [31:0] _T_2316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4252;
  reg [31:0] _T_2316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4253;
  reg [31:0] _T_2317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4254;
  reg [31:0] _T_2317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4255;
  reg [31:0] _T_2318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4256;
  reg [31:0] _T_2318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4257;
  reg [31:0] _T_2319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4258;
  reg [31:0] _T_2319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4259;
  reg [31:0] _T_2320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4260;
  reg [31:0] _T_2320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4261;
  reg [31:0] _T_2321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4262;
  reg [31:0] _T_2321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4263;
  reg [31:0] _T_2322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4264;
  reg [31:0] _T_2322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4265;
  reg [31:0] _T_2323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4266;
  reg [31:0] _T_2323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4267;
  reg [31:0] _T_2324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4268;
  reg [31:0] _T_2324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4269;
  reg [31:0] _T_2325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4270;
  reg [31:0] _T_2325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4271;
  reg [31:0] _T_2326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4272;
  reg [31:0] _T_2326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4273;
  reg [31:0] _T_2327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4274;
  reg [31:0] _T_2327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4275;
  reg [31:0] _T_2328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4276;
  reg [31:0] _T_2328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4277;
  reg [31:0] _T_2329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4278;
  reg [31:0] _T_2329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4279;
  reg [31:0] _T_2330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4280;
  reg [31:0] _T_2330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4281;
  reg [31:0] _T_2331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4282;
  reg [31:0] _T_2331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4283;
  reg [31:0] _T_2332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4284;
  reg [31:0] _T_2332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4285;
  reg [31:0] _T_2333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4286;
  reg [31:0] _T_2333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4287;
  reg [31:0] _T_2334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4288;
  reg [31:0] _T_2334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4289;
  reg [31:0] _T_2335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4290;
  reg [31:0] _T_2335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4291;
  reg [31:0] _T_2336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4292;
  reg [31:0] _T_2336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4293;
  reg [31:0] _T_2337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4294;
  reg [31:0] _T_2337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4295;
  reg [31:0] _T_2338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4296;
  reg [31:0] _T_2338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4297;
  reg [31:0] _T_2339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4298;
  reg [31:0] _T_2339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4299;
  reg [31:0] _T_2340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4300;
  reg [31:0] _T_2340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4301;
  reg [31:0] _T_2341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4302;
  reg [31:0] _T_2341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4303;
  reg [31:0] _T_2342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4304;
  reg [31:0] _T_2342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4305;
  reg [31:0] _T_2343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4306;
  reg [31:0] _T_2343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4307;
  reg [31:0] _T_2344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4308;
  reg [31:0] _T_2344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4309;
  reg [31:0] _T_2345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4310;
  reg [31:0] _T_2345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4311;
  reg [31:0] _T_2346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4312;
  reg [31:0] _T_2346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4313;
  reg [31:0] _T_2347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4314;
  reg [31:0] _T_2347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4315;
  reg [31:0] _T_2348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4316;
  reg [31:0] _T_2348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4317;
  reg [31:0] _T_2349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4318;
  reg [31:0] _T_2349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4319;
  reg [31:0] _T_2350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4320;
  reg [31:0] _T_2350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4321;
  reg [31:0] _T_2351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4322;
  reg [31:0] _T_2351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4323;
  reg [31:0] _T_2352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4324;
  reg [31:0] _T_2352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4325;
  reg [31:0] _T_2353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4326;
  reg [31:0] _T_2353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4327;
  reg [31:0] _T_2354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4328;
  reg [31:0] _T_2354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4329;
  reg [31:0] _T_2355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4330;
  reg [31:0] _T_2355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4331;
  reg [31:0] _T_2356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4332;
  reg [31:0] _T_2356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4333;
  reg [31:0] _T_2357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4334;
  reg [31:0] _T_2357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4335;
  reg [31:0] _T_2358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4336;
  reg [31:0] _T_2358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4337;
  reg [31:0] _T_2359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4338;
  reg [31:0] _T_2359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4339;
  reg [31:0] _T_2360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4340;
  reg [31:0] _T_2360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4341;
  reg [31:0] _T_2361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4342;
  reg [31:0] _T_2361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4343;
  reg [31:0] _T_2362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4344;
  reg [31:0] _T_2362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4345;
  reg [31:0] _T_2363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4346;
  reg [31:0] _T_2363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4347;
  reg [31:0] _T_2364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4348;
  reg [31:0] _T_2364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4349;
  reg [31:0] _T_2365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4350;
  reg [31:0] _T_2365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4351;
  reg [31:0] _T_2366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4352;
  reg [31:0] _T_2366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4353;
  reg [31:0] _T_2367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4354;
  reg [31:0] _T_2367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4355;
  reg [31:0] _T_2368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4356;
  reg [31:0] _T_2368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4357;
  reg [31:0] _T_2369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4358;
  reg [31:0] _T_2369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4359;
  reg [31:0] _T_2370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4360;
  reg [31:0] _T_2370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4361;
  reg [31:0] _T_2371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4362;
  reg [31:0] _T_2371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4363;
  reg [31:0] _T_2372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4364;
  reg [31:0] _T_2372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4365;
  reg [31:0] _T_2373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4366;
  reg [31:0] _T_2373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4367;
  reg [31:0] _T_2374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4368;
  reg [31:0] _T_2374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4369;
  reg [31:0] _T_2375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4370;
  reg [31:0] _T_2375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4371;
  reg [31:0] _T_2376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4372;
  reg [31:0] _T_2376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4373;
  reg [31:0] _T_2377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4374;
  reg [31:0] _T_2377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4375;
  reg [31:0] _T_2378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4376;
  reg [31:0] _T_2378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4377;
  reg [31:0] _T_2379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4378;
  reg [31:0] _T_2379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4379;
  reg [31:0] _T_2380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4380;
  reg [31:0] _T_2380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4381;
  reg [31:0] _T_2381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4382;
  reg [31:0] _T_2381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4383;
  reg [31:0] _T_2382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4384;
  reg [31:0] _T_2382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4385;
  reg [31:0] _T_2383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4386;
  reg [31:0] _T_2383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4387;
  reg [31:0] _T_2384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4388;
  reg [31:0] _T_2384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4389;
  reg [31:0] _T_2385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4390;
  reg [31:0] _T_2385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4391;
  reg [31:0] _T_2386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4392;
  reg [31:0] _T_2386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4393;
  reg [31:0] _T_2387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4394;
  reg [31:0] _T_2387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4395;
  reg [31:0] _T_2388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4396;
  reg [31:0] _T_2388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4397;
  reg [31:0] _T_2389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4398;
  reg [31:0] _T_2389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4399;
  reg [31:0] _T_2390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4400;
  reg [31:0] _T_2390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4401;
  reg [31:0] _T_2391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4402;
  reg [31:0] _T_2391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4403;
  reg [31:0] _T_2392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4404;
  reg [31:0] _T_2392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4405;
  reg [31:0] _T_2393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4406;
  reg [31:0] _T_2393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4407;
  reg [31:0] _T_2394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4408;
  reg [31:0] _T_2394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4409;
  reg [31:0] _T_2395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4410;
  reg [31:0] _T_2395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4411;
  reg [31:0] _T_2396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4412;
  reg [31:0] _T_2396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4413;
  reg [31:0] _T_2397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4414;
  reg [31:0] _T_2397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4415;
  reg [31:0] _T_2398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4416;
  reg [31:0] _T_2398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4417;
  reg [31:0] _T_2399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4418;
  reg [31:0] _T_2399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4419;
  reg [31:0] _T_2400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4420;
  reg [31:0] _T_2400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4421;
  reg [31:0] _T_2401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4422;
  reg [31:0] _T_2401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4423;
  reg [31:0] _T_2402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4424;
  reg [31:0] _T_2402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4425;
  reg [31:0] _T_2403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4426;
  reg [31:0] _T_2403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4427;
  reg [31:0] _T_2404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4428;
  reg [31:0] _T_2404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4429;
  reg [31:0] _T_2405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4430;
  reg [31:0] _T_2405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4431;
  reg [31:0] _T_2406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4432;
  reg [31:0] _T_2406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4433;
  reg [31:0] _T_2407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4434;
  reg [31:0] _T_2407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4435;
  reg [31:0] _T_2408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4436;
  reg [31:0] _T_2408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4437;
  reg [31:0] _T_2409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4438;
  reg [31:0] _T_2409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4439;
  reg [31:0] _T_2410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4440;
  reg [31:0] _T_2410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4441;
  reg [31:0] _T_2411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4442;
  reg [31:0] _T_2411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4443;
  reg [31:0] _T_2412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4444;
  reg [31:0] _T_2412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4445;
  reg [31:0] _T_2413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4446;
  reg [31:0] _T_2413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4447;
  reg [31:0] _T_2414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4448;
  reg [31:0] _T_2414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4449;
  reg [31:0] _T_2415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4450;
  reg [31:0] _T_2415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4451;
  reg [31:0] _T_2416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4452;
  reg [31:0] _T_2416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4453;
  reg [31:0] _T_2417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4454;
  reg [31:0] _T_2417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4455;
  reg [31:0] _T_2418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4456;
  reg [31:0] _T_2418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4457;
  reg [31:0] _T_2419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4458;
  reg [31:0] _T_2419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4459;
  reg [31:0] _T_2420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4460;
  reg [31:0] _T_2420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4461;
  reg [31:0] _T_2421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4462;
  reg [31:0] _T_2421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4463;
  reg [31:0] _T_2422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4464;
  reg [31:0] _T_2422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4465;
  reg [31:0] _T_2423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4466;
  reg [31:0] _T_2423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4467;
  reg [31:0] _T_2424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4468;
  reg [31:0] _T_2424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4469;
  reg [31:0] _T_2425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4470;
  reg [31:0] _T_2425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4471;
  reg [31:0] _T_2426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4472;
  reg [31:0] _T_2426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4473;
  reg [31:0] _T_2427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4474;
  reg [31:0] _T_2427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4475;
  reg [31:0] _T_2428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4476;
  reg [31:0] _T_2428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4477;
  reg [31:0] _T_2429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4478;
  reg [31:0] _T_2429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4479;
  reg [31:0] _T_2430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4480;
  reg [31:0] _T_2430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4481;
  reg [31:0] _T_2431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4482;
  reg [31:0] _T_2431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4483;
  reg [31:0] _T_2432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4484;
  reg [31:0] _T_2432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4485;
  reg [31:0] _T_2433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4486;
  reg [31:0] _T_2433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4487;
  reg [31:0] _T_2434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4488;
  reg [31:0] _T_2434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4489;
  reg [31:0] _T_2435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4490;
  reg [31:0] _T_2435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4491;
  reg [31:0] _T_2436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4492;
  reg [31:0] _T_2436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4493;
  reg [31:0] _T_2437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4494;
  reg [31:0] _T_2437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4495;
  reg [31:0] _T_2438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4496;
  reg [31:0] _T_2438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4497;
  reg [31:0] _T_2439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4498;
  reg [31:0] _T_2439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4499;
  reg [31:0] _T_2440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4500;
  reg [31:0] _T_2440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4501;
  reg [31:0] _T_2441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4502;
  reg [31:0] _T_2441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4503;
  reg [31:0] _T_2442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4504;
  reg [31:0] _T_2442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4505;
  reg [31:0] _T_2443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4506;
  reg [31:0] _T_2443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4507;
  reg [31:0] _T_2444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4508;
  reg [31:0] _T_2444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4509;
  reg [31:0] _T_2445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4510;
  reg [31:0] _T_2445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4511;
  reg [31:0] _T_2446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4512;
  reg [31:0] _T_2446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4513;
  reg [31:0] _T_2447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4514;
  reg [31:0] _T_2447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4515;
  reg [31:0] _T_2448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4516;
  reg [31:0] _T_2448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4517;
  reg [31:0] _T_2449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4518;
  reg [31:0] _T_2449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4519;
  reg [31:0] _T_2450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4520;
  reg [31:0] _T_2450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4521;
  reg [31:0] _T_2451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4522;
  reg [31:0] _T_2451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4523;
  reg [31:0] _T_2452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4524;
  reg [31:0] _T_2452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4525;
  reg [31:0] _T_2453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4526;
  reg [31:0] _T_2453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4527;
  reg [31:0] _T_2454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4528;
  reg [31:0] _T_2454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4529;
  reg [31:0] _T_2455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4530;
  reg [31:0] _T_2455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4531;
  reg [31:0] _T_2456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4532;
  reg [31:0] _T_2456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4533;
  reg [31:0] _T_2457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4534;
  reg [31:0] _T_2457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4535;
  reg [31:0] _T_2458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4536;
  reg [31:0] _T_2458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4537;
  reg [31:0] _T_2459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4538;
  reg [31:0] _T_2459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4539;
  reg [31:0] _T_2460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4540;
  reg [31:0] _T_2460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4541;
  reg [31:0] _T_2461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4542;
  reg [31:0] _T_2461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4543;
  reg [31:0] _T_2462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4544;
  reg [31:0] _T_2462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4545;
  reg [31:0] _T_2463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4546;
  reg [31:0] _T_2463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4547;
  reg [31:0] _T_2464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4548;
  reg [31:0] _T_2464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4549;
  reg [31:0] _T_2465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4550;
  reg [31:0] _T_2465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4551;
  reg [31:0] _T_2466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4552;
  reg [31:0] _T_2466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4553;
  reg [31:0] _T_2467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4554;
  reg [31:0] _T_2467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4555;
  reg [31:0] _T_2468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4556;
  reg [31:0] _T_2468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4557;
  reg [31:0] _T_2469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4558;
  reg [31:0] _T_2469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4559;
  reg [31:0] _T_2470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4560;
  reg [31:0] _T_2470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4561;
  reg [31:0] _T_2471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4562;
  reg [31:0] _T_2471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4563;
  reg [31:0] _T_2472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4564;
  reg [31:0] _T_2472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4565;
  reg [31:0] _T_2473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4566;
  reg [31:0] _T_2473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4567;
  reg [31:0] _T_2474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4568;
  reg [31:0] _T_2474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4569;
  reg [31:0] _T_2475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4570;
  reg [31:0] _T_2475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4571;
  reg [31:0] _T_2476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4572;
  reg [31:0] _T_2476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4573;
  reg [31:0] _T_2477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4574;
  reg [31:0] _T_2477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4575;
  reg [31:0] _T_2478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4576;
  reg [31:0] _T_2478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4577;
  reg [31:0] _T_2479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4578;
  reg [31:0] _T_2479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4579;
  reg [31:0] _T_2480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4580;
  reg [31:0] _T_2480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4581;
  reg [31:0] _T_2481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4582;
  reg [31:0] _T_2481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4583;
  reg [31:0] _T_2482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4584;
  reg [31:0] _T_2482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4585;
  reg [31:0] _T_2483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4586;
  reg [31:0] _T_2483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4587;
  reg [31:0] _T_2484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4588;
  reg [31:0] _T_2484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4589;
  reg [31:0] _T_2485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4590;
  reg [31:0] _T_2485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4591;
  reg [31:0] _T_2486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4592;
  reg [31:0] _T_2486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4593;
  reg [31:0] _T_2487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4594;
  reg [31:0] _T_2487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4595;
  reg [31:0] _T_2488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4596;
  reg [31:0] _T_2488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4597;
  reg [31:0] _T_2489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4598;
  reg [31:0] _T_2489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4599;
  reg [31:0] _T_2490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4600;
  reg [31:0] _T_2490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4601;
  reg [31:0] _T_2491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4602;
  reg [31:0] _T_2491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4603;
  reg [31:0] _T_2492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4604;
  reg [31:0] _T_2492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4605;
  reg [31:0] _T_2493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4606;
  reg [31:0] _T_2493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4607;
  reg [31:0] _T_2494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4608;
  reg [31:0] _T_2494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4609;
  reg [31:0] _T_2495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4610;
  reg [31:0] _T_2495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4611;
  reg [31:0] _T_2496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4612;
  reg [31:0] _T_2496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4613;
  reg [31:0] _T_2497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4614;
  reg [31:0] _T_2497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4615;
  reg [31:0] _T_2498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4616;
  reg [31:0] _T_2498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4617;
  reg [31:0] _T_2499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4618;
  reg [31:0] _T_2499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4619;
  reg [31:0] _T_2500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4620;
  reg [31:0] _T_2500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4621;
  reg [31:0] _T_2501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4622;
  reg [31:0] _T_2501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4623;
  reg [31:0] _T_2502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4624;
  reg [31:0] _T_2502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4625;
  reg [31:0] _T_2503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4626;
  reg [31:0] _T_2503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4627;
  reg [31:0] _T_2504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4628;
  reg [31:0] _T_2504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4629;
  reg [31:0] _T_2505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4630;
  reg [31:0] _T_2505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4631;
  reg [31:0] _T_2506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4632;
  reg [31:0] _T_2506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4633;
  reg [31:0] _T_2507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4634;
  reg [31:0] _T_2507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4635;
  reg [31:0] _T_2508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4636;
  reg [31:0] _T_2508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4637;
  reg [31:0] _T_2509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4638;
  reg [31:0] _T_2509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4639;
  reg [31:0] _T_2510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4640;
  reg [31:0] _T_2510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4641;
  reg [31:0] _T_2511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4642;
  reg [31:0] _T_2511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4643;
  reg [31:0] _T_2512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4644;
  reg [31:0] _T_2512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4645;
  reg [31:0] _T_2513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4646;
  reg [31:0] _T_2513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4647;
  reg [31:0] _T_2514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4648;
  reg [31:0] _T_2514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4649;
  reg [31:0] _T_2515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4650;
  reg [31:0] _T_2515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4651;
  reg [31:0] _T_2516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4652;
  reg [31:0] _T_2516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4653;
  reg [31:0] _T_2517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4654;
  reg [31:0] _T_2517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4655;
  reg [31:0] _T_2518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4656;
  reg [31:0] _T_2518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4657;
  reg [31:0] _T_2519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4658;
  reg [31:0] _T_2519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4659;
  reg [31:0] _T_2520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4660;
  reg [31:0] _T_2520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4661;
  reg [31:0] _T_2521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4662;
  reg [31:0] _T_2521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4663;
  reg [31:0] _T_2522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4664;
  reg [31:0] _T_2522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4665;
  reg [31:0] _T_2523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4666;
  reg [31:0] _T_2523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4667;
  reg [31:0] _T_2524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4668;
  reg [31:0] _T_2524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4669;
  reg [31:0] _T_2525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4670;
  reg [31:0] _T_2525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4671;
  reg [31:0] _T_2526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4672;
  reg [31:0] _T_2526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4673;
  reg [31:0] _T_2527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4674;
  reg [31:0] _T_2527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4675;
  reg [31:0] _T_2528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4676;
  reg [31:0] _T_2528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4677;
  reg [31:0] _T_2529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4678;
  reg [31:0] _T_2529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4679;
  reg [31:0] _T_2530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4680;
  reg [31:0] _T_2530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4681;
  reg [31:0] _T_2531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4682;
  reg [31:0] _T_2531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4683;
  reg [31:0] _T_2532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4684;
  reg [31:0] _T_2532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4685;
  reg [31:0] _T_2533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4686;
  reg [31:0] _T_2533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4687;
  reg [31:0] _T_2534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4688;
  reg [31:0] _T_2534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4689;
  reg [31:0] _T_2535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4690;
  reg [31:0] _T_2535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4691;
  reg [31:0] _T_2536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4692;
  reg [31:0] _T_2536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4693;
  reg [31:0] _T_2537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4694;
  reg [31:0] _T_2537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4695;
  reg [31:0] _T_2538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4696;
  reg [31:0] _T_2538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4697;
  reg [31:0] _T_2539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4698;
  reg [31:0] _T_2539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4699;
  reg [31:0] _T_2540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4700;
  reg [31:0] _T_2540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4701;
  reg [31:0] _T_2541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4702;
  reg [31:0] _T_2541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4703;
  reg [31:0] _T_2542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4704;
  reg [31:0] _T_2542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4705;
  reg [31:0] _T_2543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4706;
  reg [31:0] _T_2543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4707;
  reg [31:0] _T_2544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4708;
  reg [31:0] _T_2544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4709;
  reg [31:0] _T_2545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4710;
  reg [31:0] _T_2545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4711;
  reg [31:0] _T_2546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4712;
  reg [31:0] _T_2546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4713;
  reg [31:0] _T_2547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4714;
  reg [31:0] _T_2547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4715;
  reg [31:0] _T_2548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4716;
  reg [31:0] _T_2548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4717;
  reg [31:0] _T_2549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4718;
  reg [31:0] _T_2549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4719;
  reg [31:0] _T_2550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4720;
  reg [31:0] _T_2550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4721;
  reg [31:0] _T_2551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4722;
  reg [31:0] _T_2551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4723;
  reg [31:0] _T_2552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4724;
  reg [31:0] _T_2552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4725;
  reg [31:0] _T_2553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4726;
  reg [31:0] _T_2553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4727;
  reg [31:0] _T_2554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4728;
  reg [31:0] _T_2554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4729;
  reg [31:0] _T_2555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4730;
  reg [31:0] _T_2555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4731;
  reg [31:0] _T_2556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4732;
  reg [31:0] _T_2556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4733;
  reg [31:0] _T_2557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4734;
  reg [31:0] _T_2557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4735;
  reg [31:0] _T_2558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4736;
  reg [31:0] _T_2558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4737;
  reg [31:0] _T_2559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4738;
  reg [31:0] _T_2559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4739;
  reg [31:0] _T_2560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4740;
  reg [31:0] _T_2560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4741;
  reg [31:0] _T_2561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4742;
  reg [31:0] _T_2561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4743;
  reg [31:0] _T_2562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4744;
  reg [31:0] _T_2562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4745;
  reg [31:0] _T_2563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4746;
  reg [31:0] _T_2563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4747;
  reg [31:0] _T_2564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4748;
  reg [31:0] _T_2564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4749;
  reg [31:0] _T_2565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4750;
  reg [31:0] _T_2565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4751;
  reg [31:0] _T_2566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4752;
  reg [31:0] _T_2566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4753;
  reg [31:0] _T_2567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4754;
  reg [31:0] _T_2567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4755;
  reg [31:0] _T_2568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4756;
  reg [31:0] _T_2568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4757;
  reg [31:0] _T_2569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4758;
  reg [31:0] _T_2569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4759;
  reg [31:0] _T_2570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4760;
  reg [31:0] _T_2570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4761;
  reg [31:0] _T_2571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4762;
  reg [31:0] _T_2571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4763;
  reg [31:0] _T_2572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4764;
  reg [31:0] _T_2572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4765;
  reg [31:0] _T_2573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4766;
  reg [31:0] _T_2573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4767;
  reg [31:0] _T_2574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4768;
  reg [31:0] _T_2574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4769;
  reg [31:0] _T_2575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4770;
  reg [31:0] _T_2575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4771;
  reg [31:0] _T_2576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4772;
  reg [31:0] _T_2576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4773;
  reg [31:0] _T_2577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4774;
  reg [31:0] _T_2577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4775;
  reg [31:0] _T_2578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4776;
  reg [31:0] _T_2578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4777;
  reg [31:0] _T_2579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4778;
  reg [31:0] _T_2579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4779;
  reg [31:0] _T_2580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4780;
  reg [31:0] _T_2580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4781;
  reg [31:0] _T_2581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4782;
  reg [31:0] _T_2581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4783;
  reg [31:0] _T_2582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4784;
  reg [31:0] _T_2582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4785;
  reg [31:0] _T_2583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4786;
  reg [31:0] _T_2583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4787;
  reg [31:0] _T_2584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4788;
  reg [31:0] _T_2584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4789;
  reg [31:0] _T_2585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4790;
  reg [31:0] _T_2585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4791;
  reg [31:0] _T_2586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4792;
  reg [31:0] _T_2586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4793;
  reg [31:0] _T_2587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4794;
  reg [31:0] _T_2587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4795;
  reg [31:0] _T_2588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4796;
  reg [31:0] _T_2588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4797;
  reg [31:0] _T_2589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4798;
  reg [31:0] _T_2589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4799;
  reg [31:0] _T_2590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4800;
  reg [31:0] _T_2590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4801;
  reg [31:0] _T_2591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4802;
  reg [31:0] _T_2591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4803;
  reg [31:0] _T_2592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4804;
  reg [31:0] _T_2592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4805;
  reg [31:0] _T_2593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4806;
  reg [31:0] _T_2593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4807;
  reg [31:0] _T_2594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4808;
  reg [31:0] _T_2594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4809;
  reg [31:0] _T_2595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4810;
  reg [31:0] _T_2595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4811;
  reg [31:0] _T_2596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4812;
  reg [31:0] _T_2596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4813;
  reg [31:0] _T_2597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4814;
  reg [31:0] _T_2597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4815;
  reg [31:0] _T_2598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4816;
  reg [31:0] _T_2598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4817;
  reg [31:0] _T_2599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4818;
  reg [31:0] _T_2599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4819;
  reg [31:0] _T_2600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4820;
  reg [31:0] _T_2600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4821;
  reg [31:0] _T_2601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4822;
  reg [31:0] _T_2601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4823;
  reg [31:0] _T_2602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4824;
  reg [31:0] _T_2602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4825;
  reg [31:0] _T_2603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4826;
  reg [31:0] _T_2603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4827;
  reg [31:0] _T_2604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4828;
  reg [31:0] _T_2604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4829;
  reg [31:0] _T_2605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4830;
  reg [31:0] _T_2605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4831;
  reg [31:0] _T_2606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4832;
  reg [31:0] _T_2606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4833;
  reg [31:0] _T_2607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4834;
  reg [31:0] _T_2607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4835;
  reg [31:0] _T_2608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4836;
  reg [31:0] _T_2608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4837;
  reg [31:0] _T_2609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4838;
  reg [31:0] _T_2609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4839;
  reg [31:0] _T_2610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4840;
  reg [31:0] _T_2610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4841;
  reg [31:0] _T_2611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4842;
  reg [31:0] _T_2611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4843;
  reg [31:0] _T_2612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4844;
  reg [31:0] _T_2612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4845;
  reg [31:0] _T_2613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4846;
  reg [31:0] _T_2613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4847;
  reg [31:0] _T_2614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4848;
  reg [31:0] _T_2614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4849;
  reg [31:0] _T_2615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4850;
  reg [31:0] _T_2615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4851;
  reg [31:0] _T_2616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4852;
  reg [31:0] _T_2616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4853;
  reg [31:0] _T_2617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4854;
  reg [31:0] _T_2617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4855;
  reg [31:0] _T_2618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4856;
  reg [31:0] _T_2618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4857;
  reg [31:0] _T_2619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4858;
  reg [31:0] _T_2619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4859;
  reg [31:0] _T_2620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4860;
  reg [31:0] _T_2620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4861;
  reg [31:0] _T_2621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4862;
  reg [31:0] _T_2621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4863;
  reg [31:0] _T_2622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4864;
  reg [31:0] _T_2622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4865;
  reg [31:0] _T_2623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4866;
  reg [31:0] _T_2623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4867;
  reg [31:0] _T_2624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4868;
  reg [31:0] _T_2624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4869;
  reg [31:0] _T_2625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4870;
  reg [31:0] _T_2625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4871;
  reg [31:0] _T_2626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4872;
  reg [31:0] _T_2626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4873;
  reg [31:0] _T_2627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4874;
  reg [31:0] _T_2627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4875;
  reg [31:0] _T_2628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4876;
  reg [31:0] _T_2628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4877;
  reg [31:0] _T_2629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4878;
  reg [31:0] _T_2629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4879;
  reg [31:0] _T_2630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4880;
  reg [31:0] _T_2630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4881;
  reg [31:0] _T_2631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4882;
  reg [31:0] _T_2631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4883;
  reg [31:0] _T_2632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4884;
  reg [31:0] _T_2632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4885;
  reg [31:0] _T_2633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4886;
  reg [31:0] _T_2633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4887;
  reg [31:0] _T_2634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4888;
  reg [31:0] _T_2634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4889;
  reg [31:0] _T_2635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4890;
  reg [31:0] _T_2635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4891;
  reg [31:0] _T_2636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4892;
  reg [31:0] _T_2636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4893;
  reg [31:0] _T_2637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4894;
  reg [31:0] _T_2637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4895;
  reg [31:0] _T_2638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4896;
  reg [31:0] _T_2638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4897;
  reg [31:0] _T_2639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4898;
  reg [31:0] _T_2639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4899;
  reg [31:0] _T_2640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4900;
  reg [31:0] _T_2640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4901;
  reg [31:0] _T_2641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4902;
  reg [31:0] _T_2641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4903;
  reg [31:0] _T_2642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4904;
  reg [31:0] _T_2642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4905;
  reg [31:0] _T_2643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4906;
  reg [31:0] _T_2643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4907;
  reg [31:0] _T_2644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4908;
  reg [31:0] _T_2644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4909;
  reg [31:0] _T_2645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4910;
  reg [31:0] _T_2645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4911;
  reg [31:0] _T_2646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4912;
  reg [31:0] _T_2646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4913;
  reg [31:0] _T_2647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4914;
  reg [31:0] _T_2647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4915;
  reg [31:0] _T_2648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4916;
  reg [31:0] _T_2648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4917;
  reg [31:0] _T_2649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4918;
  reg [31:0] _T_2649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4919;
  reg [31:0] _T_2650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4920;
  reg [31:0] _T_2650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4921;
  reg [31:0] _T_2651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4922;
  reg [31:0] _T_2651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4923;
  reg [31:0] _T_2652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4924;
  reg [31:0] _T_2652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4925;
  reg [31:0] _T_2653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4926;
  reg [31:0] _T_2653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4927;
  reg [31:0] _T_2654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4928;
  reg [31:0] _T_2654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4929;
  reg [31:0] _T_2655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4930;
  reg [31:0] _T_2655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4931;
  reg [31:0] _T_2656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4932;
  reg [31:0] _T_2656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4933;
  reg [31:0] _T_2657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4934;
  reg [31:0] _T_2657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4935;
  reg [31:0] _T_2658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4936;
  reg [31:0] _T_2658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4937;
  reg [31:0] _T_2659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4938;
  reg [31:0] _T_2659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4939;
  reg [31:0] _T_2660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4940;
  reg [31:0] _T_2660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4941;
  reg [31:0] _T_2661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4942;
  reg [31:0] _T_2661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4943;
  reg [31:0] _T_2662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4944;
  reg [31:0] _T_2662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4945;
  reg [31:0] _T_2663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4946;
  reg [31:0] _T_2663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4947;
  reg [31:0] _T_2664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4948;
  reg [31:0] _T_2664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4949;
  reg [31:0] _T_2665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4950;
  reg [31:0] _T_2665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4951;
  reg [31:0] _T_2666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4952;
  reg [31:0] _T_2666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4953;
  reg [31:0] _T_2667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4954;
  reg [31:0] _T_2667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4955;
  reg [31:0] _T_2668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4956;
  reg [31:0] _T_2668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4957;
  reg [31:0] _T_2669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4958;
  reg [31:0] _T_2669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4959;
  reg [31:0] _T_2670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4960;
  reg [31:0] _T_2670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4961;
  reg [31:0] _T_2671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4962;
  reg [31:0] _T_2671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4963;
  reg [31:0] _T_2672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4964;
  reg [31:0] _T_2672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4965;
  reg [31:0] _T_2673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4966;
  reg [31:0] _T_2673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4967;
  reg [31:0] _T_2674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4968;
  reg [31:0] _T_2674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4969;
  reg [31:0] _T_2675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4970;
  reg [31:0] _T_2675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4971;
  reg [31:0] _T_2676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4972;
  reg [31:0] _T_2676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4973;
  reg [31:0] _T_2677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4974;
  reg [31:0] _T_2677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4975;
  reg [31:0] _T_2678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4976;
  reg [31:0] _T_2678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4977;
  reg [31:0] _T_2679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4978;
  reg [31:0] _T_2679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4979;
  reg [31:0] _T_2680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4980;
  reg [31:0] _T_2680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4981;
  reg [31:0] _T_2681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4982;
  reg [31:0] _T_2681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4983;
  reg [31:0] _T_2682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4984;
  reg [31:0] _T_2682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4985;
  reg [31:0] _T_2683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4986;
  reg [31:0] _T_2683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4987;
  reg [31:0] _T_2684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4988;
  reg [31:0] _T_2684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4989;
  reg [31:0] _T_2685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4990;
  reg [31:0] _T_2685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4991;
  reg [31:0] _T_2686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4992;
  reg [31:0] _T_2686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4993;
  reg [31:0] _T_2687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4994;
  reg [31:0] _T_2687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4995;
  reg [31:0] _T_2688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4996;
  reg [31:0] _T_2688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4997;
  reg [31:0] _T_2689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4998;
  reg [31:0] _T_2689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4999;
  reg [31:0] _T_2690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5000;
  reg [31:0] _T_2690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5001;
  reg [31:0] _T_2691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5002;
  reg [31:0] _T_2691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5003;
  reg [31:0] _T_2692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5004;
  reg [31:0] _T_2692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5005;
  reg [31:0] _T_2693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5006;
  reg [31:0] _T_2693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5007;
  reg [31:0] _T_2694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5008;
  reg [31:0] _T_2694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5009;
  reg [31:0] _T_2695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5010;
  reg [31:0] _T_2695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5011;
  reg [31:0] _T_2696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5012;
  reg [31:0] _T_2696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5013;
  reg [31:0] _T_2697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5014;
  reg [31:0] _T_2697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5015;
  reg [31:0] _T_2698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5016;
  reg [31:0] _T_2698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5017;
  reg [31:0] _T_2699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5018;
  reg [31:0] _T_2699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5019;
  reg [31:0] _T_2700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5020;
  reg [31:0] _T_2700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5021;
  reg [31:0] _T_2701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5022;
  reg [31:0] _T_2701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5023;
  reg [31:0] _T_2702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5024;
  reg [31:0] _T_2702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5025;
  reg [31:0] _T_2703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5026;
  reg [31:0] _T_2703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5027;
  reg [31:0] _T_2704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5028;
  reg [31:0] _T_2704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5029;
  reg [31:0] _T_2705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5030;
  reg [31:0] _T_2705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5031;
  reg [31:0] _T_2706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5032;
  reg [31:0] _T_2706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5033;
  reg [31:0] _T_2707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5034;
  reg [31:0] _T_2707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5035;
  reg [31:0] _T_2708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5036;
  reg [31:0] _T_2708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5037;
  reg [31:0] _T_2709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5038;
  reg [31:0] _T_2709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5039;
  reg [31:0] _T_2710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5040;
  reg [31:0] _T_2710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5041;
  reg [31:0] _T_2711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5042;
  reg [31:0] _T_2711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5043;
  reg [31:0] _T_2712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5044;
  reg [31:0] _T_2712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5045;
  reg [31:0] _T_2713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5046;
  reg [31:0] _T_2713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5047;
  reg [31:0] _T_2714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5048;
  reg [31:0] _T_2714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5049;
  reg [31:0] _T_2715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5050;
  reg [31:0] _T_2715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5051;
  reg [31:0] _T_2716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5052;
  reg [31:0] _T_2716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5053;
  reg [31:0] _T_2717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5054;
  reg [31:0] _T_2717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5055;
  reg [31:0] _T_2718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5056;
  reg [31:0] _T_2718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5057;
  reg [31:0] _T_2719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5058;
  reg [31:0] _T_2719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5059;
  reg [31:0] _T_2720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5060;
  reg [31:0] _T_2720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5061;
  reg [31:0] _T_2721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5062;
  reg [31:0] _T_2721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5063;
  reg [31:0] _T_2722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5064;
  reg [31:0] _T_2722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5065;
  reg [31:0] _T_2723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5066;
  reg [31:0] _T_2723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5067;
  reg [31:0] _T_2724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5068;
  reg [31:0] _T_2724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5069;
  reg [31:0] _T_2725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5070;
  reg [31:0] _T_2725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5071;
  reg [31:0] _T_2726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5072;
  reg [31:0] _T_2726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5073;
  reg [31:0] _T_2727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5074;
  reg [31:0] _T_2727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5075;
  reg [31:0] _T_2728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5076;
  reg [31:0] _T_2728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5077;
  reg [31:0] _T_2729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5078;
  reg [31:0] _T_2729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5079;
  reg [31:0] _T_2730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5080;
  reg [31:0] _T_2730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5081;
  reg [31:0] _T_2731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5082;
  reg [31:0] _T_2731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5083;
  reg [31:0] _T_2732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5084;
  reg [31:0] _T_2732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5085;
  reg [31:0] _T_2733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5086;
  reg [31:0] _T_2733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5087;
  reg [31:0] _T_2734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5088;
  reg [31:0] _T_2734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5089;
  reg [31:0] _T_2735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5090;
  reg [31:0] _T_2735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5091;
  reg [31:0] _T_2736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5092;
  reg [31:0] _T_2736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5093;
  reg [31:0] _T_2737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5094;
  reg [31:0] _T_2737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5095;
  reg [31:0] _T_2738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5096;
  reg [31:0] _T_2738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5097;
  reg [31:0] _T_2739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5098;
  reg [31:0] _T_2739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5099;
  reg [31:0] _T_2740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5100;
  reg [31:0] _T_2740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5101;
  reg [31:0] _T_2741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5102;
  reg [31:0] _T_2741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5103;
  reg [31:0] _T_2742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5104;
  reg [31:0] _T_2742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5105;
  reg [31:0] _T_2743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5106;
  reg [31:0] _T_2743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5107;
  reg [31:0] _T_2744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5108;
  reg [31:0] _T_2744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5109;
  reg [31:0] _T_2745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5110;
  reg [31:0] _T_2745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5111;
  reg [31:0] _T_2746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5112;
  reg [31:0] _T_2746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5113;
  reg [31:0] _T_2747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5114;
  reg [31:0] _T_2747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5115;
  reg [31:0] _T_2748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5116;
  reg [31:0] _T_2748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5117;
  reg [31:0] _T_2749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5118;
  reg [31:0] _T_2749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5119;
  reg [31:0] _T_2750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5120;
  reg [31:0] _T_2750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5121;
  reg [31:0] _T_2751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5122;
  reg [31:0] _T_2751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5123;
  reg [31:0] _T_2752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5124;
  reg [31:0] _T_2752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5125;
  reg [31:0] _T_2753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5126;
  reg [31:0] _T_2753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5127;
  reg [31:0] _T_2754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5128;
  reg [31:0] _T_2754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5129;
  reg [31:0] _T_2755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5130;
  reg [31:0] _T_2755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5131;
  reg [31:0] _T_2756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5132;
  reg [31:0] _T_2756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5133;
  reg [31:0] _T_2757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5134;
  reg [31:0] _T_2757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5135;
  reg [31:0] _T_2758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5136;
  reg [31:0] _T_2758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5137;
  reg [31:0] _T_2759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5138;
  reg [31:0] _T_2759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5139;
  reg [31:0] _T_2760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5140;
  reg [31:0] _T_2760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5141;
  reg [31:0] _T_2761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5142;
  reg [31:0] _T_2761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5143;
  reg [31:0] _T_2762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5144;
  reg [31:0] _T_2762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5145;
  reg [31:0] _T_2763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5146;
  reg [31:0] _T_2763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5147;
  reg [31:0] _T_2764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5148;
  reg [31:0] _T_2764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5149;
  reg [31:0] _T_2765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5150;
  reg [31:0] _T_2765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5151;
  reg [31:0] _T_2766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5152;
  reg [31:0] _T_2766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5153;
  reg [31:0] _T_2767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5154;
  reg [31:0] _T_2767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5155;
  reg [31:0] _T_2768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5156;
  reg [31:0] _T_2768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5157;
  reg [31:0] _T_2769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5158;
  reg [31:0] _T_2769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5159;
  reg [31:0] _T_2770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5160;
  reg [31:0] _T_2770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5161;
  reg [31:0] _T_2771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5162;
  reg [31:0] _T_2771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5163;
  reg [31:0] _T_2772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5164;
  reg [31:0] _T_2772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5165;
  reg [31:0] _T_2773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5166;
  reg [31:0] _T_2773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5167;
  reg [31:0] _T_2774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5168;
  reg [31:0] _T_2774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5169;
  reg [31:0] _T_2775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5170;
  reg [31:0] _T_2775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5171;
  reg [31:0] _T_2776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5172;
  reg [31:0] _T_2776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5173;
  reg [31:0] _T_2777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5174;
  reg [31:0] _T_2777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5175;
  reg [31:0] _T_2778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5176;
  reg [31:0] _T_2778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5177;
  reg [31:0] _T_2779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5178;
  reg [31:0] _T_2779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5179;
  reg [31:0] _T_2780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5180;
  reg [31:0] _T_2780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5181;
  reg [31:0] _T_2781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5182;
  reg [31:0] _T_2781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5183;
  reg [31:0] _T_2782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5184;
  reg [31:0] _T_2782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5185;
  reg [31:0] _T_2783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5186;
  reg [31:0] _T_2783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5187;
  reg [31:0] _T_2784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5188;
  reg [31:0] _T_2784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5189;
  reg [31:0] _T_2785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5190;
  reg [31:0] _T_2785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5191;
  reg [31:0] _T_2786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5192;
  reg [31:0] _T_2786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5193;
  reg [31:0] _T_2787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5194;
  reg [31:0] _T_2787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5195;
  reg [31:0] _T_2788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5196;
  reg [31:0] _T_2788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5197;
  reg [31:0] _T_2789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5198;
  reg [31:0] _T_2789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5199;
  reg [31:0] _T_2790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5200;
  reg [31:0] _T_2790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5201;
  reg [31:0] _T_2791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5202;
  reg [31:0] _T_2791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5203;
  reg [31:0] _T_2792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5204;
  reg [31:0] _T_2792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5205;
  reg [31:0] _T_2793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5206;
  reg [31:0] _T_2793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5207;
  reg [31:0] _T_2794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5208;
  reg [31:0] _T_2794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5209;
  reg [31:0] _T_2795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5210;
  reg [31:0] _T_2795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5211;
  reg [31:0] _T_2796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5212;
  reg [31:0] _T_2796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5213;
  reg [31:0] _T_2797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5214;
  reg [31:0] _T_2797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5215;
  reg [31:0] _T_2798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5216;
  reg [31:0] _T_2798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5217;
  reg [31:0] _T_2799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5218;
  reg [31:0] _T_2799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5219;
  reg [31:0] _T_2800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5220;
  reg [31:0] _T_2800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5221;
  reg [31:0] _T_2801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5222;
  reg [31:0] _T_2801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5223;
  reg [31:0] _T_2802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5224;
  reg [31:0] _T_2802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5225;
  reg [31:0] _T_2803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5226;
  reg [31:0] _T_2803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5227;
  reg [31:0] _T_2804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5228;
  reg [31:0] _T_2804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5229;
  reg [31:0] _T_2805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5230;
  reg [31:0] _T_2805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5231;
  reg [31:0] _T_2806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5232;
  reg [31:0] _T_2806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5233;
  reg [31:0] _T_2807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5234;
  reg [31:0] _T_2807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5235;
  reg [31:0] _T_2808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5236;
  reg [31:0] _T_2808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5237;
  reg [31:0] _T_2809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5238;
  reg [31:0] _T_2809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5239;
  reg [31:0] _T_2810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5240;
  reg [31:0] _T_2810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5241;
  reg [31:0] _T_2811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5242;
  reg [31:0] _T_2811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5243;
  reg [31:0] _T_2812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5244;
  reg [31:0] _T_2812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5245;
  reg [31:0] _T_2813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5246;
  reg [31:0] _T_2813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5247;
  reg [31:0] _T_2814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5248;
  reg [31:0] _T_2814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5249;
  reg [31:0] _T_2815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5250;
  reg [31:0] _T_2815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5251;
  reg [31:0] _T_2816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5252;
  reg [31:0] _T_2816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5253;
  reg [31:0] _T_2817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5254;
  reg [31:0] _T_2817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5255;
  reg [31:0] _T_2818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5256;
  reg [31:0] _T_2818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5257;
  reg [31:0] _T_2819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5258;
  reg [31:0] _T_2819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5259;
  reg [31:0] _T_2820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5260;
  reg [31:0] _T_2820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5261;
  reg [31:0] _T_2821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5262;
  reg [31:0] _T_2821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5263;
  reg [31:0] _T_2822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5264;
  reg [31:0] _T_2822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5265;
  reg [31:0] _T_2823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5266;
  reg [31:0] _T_2823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5267;
  reg [31:0] _T_2824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5268;
  reg [31:0] _T_2824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5269;
  reg [31:0] _T_2825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5270;
  reg [31:0] _T_2825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5271;
  reg [31:0] _T_2826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5272;
  reg [31:0] _T_2826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5273;
  reg [31:0] _T_2827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5274;
  reg [31:0] _T_2827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5275;
  reg [31:0] _T_2828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5276;
  reg [31:0] _T_2828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5277;
  reg [31:0] _T_2829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5278;
  reg [31:0] _T_2829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5279;
  reg [31:0] _T_2830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5280;
  reg [31:0] _T_2830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5281;
  reg [31:0] _T_2831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5282;
  reg [31:0] _T_2831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5283;
  reg [31:0] _T_2832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5284;
  reg [31:0] _T_2832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5285;
  reg [31:0] _T_2833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5286;
  reg [31:0] _T_2833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5287;
  reg [31:0] _T_2834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5288;
  reg [31:0] _T_2834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5289;
  reg [31:0] _T_2835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5290;
  reg [31:0] _T_2835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5291;
  reg [31:0] _T_2836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5292;
  reg [31:0] _T_2836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5293;
  reg [31:0] _T_2837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5294;
  reg [31:0] _T_2837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5295;
  reg [31:0] _T_2838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5296;
  reg [31:0] _T_2838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5297;
  reg [31:0] _T_2839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5298;
  reg [31:0] _T_2839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5299;
  reg [31:0] _T_2840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5300;
  reg [31:0] _T_2840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5301;
  reg [31:0] _T_2841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5302;
  reg [31:0] _T_2841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5303;
  reg [31:0] _T_2842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5304;
  reg [31:0] _T_2842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5305;
  reg [31:0] _T_2843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5306;
  reg [31:0] _T_2843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5307;
  reg [31:0] _T_2844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5308;
  reg [31:0] _T_2844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5309;
  reg [31:0] _T_2845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5310;
  reg [31:0] _T_2845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5311;
  reg [31:0] _T_2846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5312;
  reg [31:0] _T_2846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5313;
  reg [31:0] _T_2847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5314;
  reg [31:0] _T_2847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5315;
  reg [31:0] _T_2848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5316;
  reg [31:0] _T_2848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5317;
  reg [31:0] _T_2849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5318;
  reg [31:0] _T_2849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5319;
  reg [31:0] _T_2850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5320;
  reg [31:0] _T_2850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5321;
  reg [31:0] _T_2851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5322;
  reg [31:0] _T_2851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5323;
  reg [31:0] _T_2852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5324;
  reg [31:0] _T_2852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5325;
  reg [31:0] _T_2853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5326;
  reg [31:0] _T_2853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5327;
  reg [31:0] _T_2854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5328;
  reg [31:0] _T_2854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5329;
  reg [31:0] _T_2855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5330;
  reg [31:0] _T_2855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5331;
  reg [31:0] _T_2856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5332;
  reg [31:0] _T_2856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5333;
  reg [31:0] _T_2857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5334;
  reg [31:0] _T_2857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5335;
  reg [31:0] _T_2858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5336;
  reg [31:0] _T_2858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5337;
  reg [31:0] _T_2859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5338;
  reg [31:0] _T_2859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5339;
  reg [31:0] _T_2860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5340;
  reg [31:0] _T_2860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5341;
  reg [31:0] _T_2861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5342;
  reg [31:0] _T_2861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5343;
  reg [31:0] _T_2862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5344;
  reg [31:0] _T_2862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5345;
  reg [31:0] _T_2863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5346;
  reg [31:0] _T_2863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5347;
  reg [31:0] _T_2864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5348;
  reg [31:0] _T_2864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5349;
  reg [31:0] _T_2865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5350;
  reg [31:0] _T_2865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5351;
  reg [31:0] _T_2866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5352;
  reg [31:0] _T_2866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5353;
  reg [31:0] _T_2867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5354;
  reg [31:0] _T_2867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5355;
  reg [31:0] _T_2868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5356;
  reg [31:0] _T_2868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5357;
  reg [31:0] _T_2869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5358;
  reg [31:0] _T_2869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5359;
  reg [31:0] _T_2870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5360;
  reg [31:0] _T_2870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5361;
  reg [31:0] _T_2871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5362;
  reg [31:0] _T_2871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5363;
  reg [31:0] _T_2872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5364;
  reg [31:0] _T_2872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5365;
  reg [31:0] _T_2873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5366;
  reg [31:0] _T_2873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5367;
  reg [31:0] _T_2874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5368;
  reg [31:0] _T_2874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5369;
  reg [31:0] _T_2875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5370;
  reg [31:0] _T_2875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5371;
  reg [31:0] _T_2876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5372;
  reg [31:0] _T_2876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5373;
  reg [31:0] _T_2877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5374;
  reg [31:0] _T_2877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5375;
  reg [31:0] _T_2878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5376;
  reg [31:0] _T_2878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5377;
  reg [31:0] _T_2879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5378;
  reg [31:0] _T_2879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5379;
  reg [31:0] _T_2880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5380;
  reg [31:0] _T_2880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5381;
  reg [31:0] _T_2881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5382;
  reg [31:0] _T_2881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5383;
  reg [31:0] _T_2882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5384;
  reg [31:0] _T_2882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5385;
  reg [31:0] _T_2883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5386;
  reg [31:0] _T_2883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5387;
  reg [31:0] _T_2884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5388;
  reg [31:0] _T_2884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5389;
  reg [31:0] _T_2885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5390;
  reg [31:0] _T_2885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5391;
  reg [31:0] _T_2886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5392;
  reg [31:0] _T_2886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5393;
  reg [31:0] _T_2887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5394;
  reg [31:0] _T_2887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5395;
  reg [31:0] _T_2888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5396;
  reg [31:0] _T_2888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5397;
  reg [31:0] _T_2889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5398;
  reg [31:0] _T_2889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5399;
  reg [31:0] _T_2890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5400;
  reg [31:0] _T_2890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5401;
  reg [31:0] _T_2891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5402;
  reg [31:0] _T_2891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5403;
  reg [31:0] _T_2892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5404;
  reg [31:0] _T_2892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5405;
  reg [31:0] _T_2893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5406;
  reg [31:0] _T_2893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5407;
  reg [31:0] _T_2894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5408;
  reg [31:0] _T_2894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5409;
  reg [31:0] _T_2895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5410;
  reg [31:0] _T_2895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5411;
  reg [31:0] _T_2896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5412;
  reg [31:0] _T_2896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5413;
  reg [31:0] _T_2897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5414;
  reg [31:0] _T_2897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5415;
  reg [31:0] _T_2898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5416;
  reg [31:0] _T_2898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5417;
  reg [31:0] _T_2899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5418;
  reg [31:0] _T_2899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5419;
  reg [31:0] _T_2900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5420;
  reg [31:0] _T_2900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5421;
  reg [31:0] _T_2901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5422;
  reg [31:0] _T_2901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5423;
  reg [31:0] _T_2902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5424;
  reg [31:0] _T_2902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5425;
  reg [31:0] _T_2903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5426;
  reg [31:0] _T_2903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5427;
  reg [31:0] _T_2904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5428;
  reg [31:0] _T_2904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5429;
  reg [31:0] _T_2905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5430;
  reg [31:0] _T_2905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5431;
  reg [31:0] _T_2906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5432;
  reg [31:0] _T_2906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5433;
  reg [31:0] _T_2907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5434;
  reg [31:0] _T_2907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5435;
  reg [31:0] _T_2908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5436;
  reg [31:0] _T_2908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5437;
  reg [31:0] _T_2909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5438;
  reg [31:0] _T_2909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5439;
  reg [31:0] _T_2910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5440;
  reg [31:0] _T_2910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5441;
  reg [31:0] _T_2911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5442;
  reg [31:0] _T_2911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5443;
  reg [31:0] _T_2912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5444;
  reg [31:0] _T_2912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5445;
  reg [31:0] _T_2913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5446;
  reg [31:0] _T_2913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5447;
  reg [31:0] _T_2914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5448;
  reg [31:0] _T_2914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5449;
  reg [31:0] _T_2915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5450;
  reg [31:0] _T_2915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5451;
  reg [31:0] _T_2916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5452;
  reg [31:0] _T_2916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5453;
  reg [31:0] _T_2917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5454;
  reg [31:0] _T_2917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5455;
  reg [31:0] _T_2918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5456;
  reg [31:0] _T_2918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5457;
  reg [31:0] _T_2919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5458;
  reg [31:0] _T_2919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5459;
  reg [31:0] _T_2920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5460;
  reg [31:0] _T_2920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5461;
  reg [31:0] _T_2921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5462;
  reg [31:0] _T_2921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5463;
  reg [31:0] _T_2922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5464;
  reg [31:0] _T_2922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5465;
  reg [31:0] _T_2923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5466;
  reg [31:0] _T_2923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5467;
  reg [31:0] _T_2924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5468;
  reg [31:0] _T_2924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5469;
  reg [31:0] _T_2925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5470;
  reg [31:0] _T_2925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5471;
  reg [31:0] _T_2926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5472;
  reg [31:0] _T_2926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5473;
  reg [31:0] _T_2927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5474;
  reg [31:0] _T_2927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5475;
  reg [31:0] _T_2928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5476;
  reg [31:0] _T_2928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5477;
  reg [31:0] _T_2929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5478;
  reg [31:0] _T_2929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5479;
  reg [31:0] _T_2930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5480;
  reg [31:0] _T_2930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5481;
  reg [31:0] _T_2931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5482;
  reg [31:0] _T_2931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5483;
  reg [31:0] _T_2932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5484;
  reg [31:0] _T_2932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5485;
  reg [31:0] _T_2933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5486;
  reg [31:0] _T_2933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5487;
  reg [31:0] _T_2934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5488;
  reg [31:0] _T_2934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5489;
  reg [31:0] _T_2935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5490;
  reg [31:0] _T_2935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5491;
  reg [31:0] _T_2936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5492;
  reg [31:0] _T_2936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5493;
  reg [31:0] _T_2937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5494;
  reg [31:0] _T_2937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5495;
  reg [31:0] _T_2938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5496;
  reg [31:0] _T_2938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5497;
  reg [31:0] _T_2939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5498;
  reg [31:0] _T_2939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5499;
  reg [31:0] _T_2940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5500;
  reg [31:0] _T_2940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5501;
  reg [31:0] _T_2941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5502;
  reg [31:0] _T_2941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5503;
  reg [31:0] _T_2942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5504;
  reg [31:0] _T_2942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5505;
  reg [31:0] _T_2943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5506;
  reg [31:0] _T_2943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5507;
  reg [31:0] _T_2944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5508;
  reg [31:0] _T_2944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5509;
  reg [31:0] _T_2945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5510;
  reg [31:0] _T_2945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5511;
  reg [31:0] _T_2946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5512;
  reg [31:0] _T_2946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5513;
  reg [31:0] _T_2947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5514;
  reg [31:0] _T_2947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5515;
  reg [31:0] _T_2948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5516;
  reg [31:0] _T_2948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5517;
  reg [31:0] _T_2949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5518;
  reg [31:0] _T_2949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5519;
  reg [31:0] _T_2950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5520;
  reg [31:0] _T_2950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5521;
  reg [31:0] _T_2951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5522;
  reg [31:0] _T_2951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5523;
  reg [31:0] _T_2952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5524;
  reg [31:0] _T_2952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5525;
  reg [31:0] _T_2953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5526;
  reg [31:0] _T_2953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5527;
  reg [31:0] _T_2954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5528;
  reg [31:0] _T_2954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5529;
  reg [31:0] _T_2955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5530;
  reg [31:0] _T_2955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5531;
  reg [31:0] _T_2956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5532;
  reg [31:0] _T_2956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5533;
  reg [31:0] _T_2957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5534;
  reg [31:0] _T_2957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5535;
  reg [31:0] _T_2958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5536;
  reg [31:0] _T_2958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5537;
  reg [31:0] _T_2959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5538;
  reg [31:0] _T_2959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5539;
  reg [31:0] _T_2960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5540;
  reg [31:0] _T_2960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5541;
  reg [31:0] _T_2961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5542;
  reg [31:0] _T_2961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5543;
  reg [31:0] _T_2962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5544;
  reg [31:0] _T_2962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5545;
  reg [31:0] _T_2963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5546;
  reg [31:0] _T_2963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5547;
  reg [31:0] _T_2964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5548;
  reg [31:0] _T_2964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5549;
  reg [31:0] _T_2965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5550;
  reg [31:0] _T_2965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5551;
  reg [31:0] _T_2966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5552;
  reg [31:0] _T_2966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5553;
  reg [31:0] _T_2967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5554;
  reg [31:0] _T_2967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5555;
  reg [31:0] _T_2968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5556;
  reg [31:0] _T_2968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5557;
  reg [31:0] _T_2969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5558;
  reg [31:0] _T_2969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5559;
  reg [31:0] _T_2970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5560;
  reg [31:0] _T_2970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5561;
  reg [31:0] _T_2971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5562;
  reg [31:0] _T_2971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5563;
  reg [31:0] _T_2972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5564;
  reg [31:0] _T_2972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5565;
  reg [31:0] _T_2973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5566;
  reg [31:0] _T_2973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5567;
  reg [31:0] _T_2974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5568;
  reg [31:0] _T_2974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5569;
  reg [31:0] _T_2975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5570;
  reg [31:0] _T_2975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5571;
  reg [31:0] _T_2976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5572;
  reg [31:0] _T_2976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5573;
  reg [31:0] _T_2977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5574;
  reg [31:0] _T_2977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5575;
  reg [31:0] _T_2978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5576;
  reg [31:0] _T_2978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5577;
  reg [31:0] _T_2979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5578;
  reg [31:0] _T_2979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5579;
  reg [31:0] _T_2980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5580;
  reg [31:0] _T_2980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5581;
  reg [31:0] _T_2981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5582;
  reg [31:0] _T_2981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5583;
  reg [31:0] _T_2982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5584;
  reg [31:0] _T_2982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5585;
  reg [31:0] _T_2983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5586;
  reg [31:0] _T_2983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5587;
  reg [31:0] _T_2984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5588;
  reg [31:0] _T_2984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5589;
  reg [31:0] _T_2985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5590;
  reg [31:0] _T_2985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5591;
  reg [31:0] _T_2986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5592;
  reg [31:0] _T_2986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5593;
  reg [31:0] _T_2987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5594;
  reg [31:0] _T_2987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5595;
  reg [31:0] _T_2988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5596;
  reg [31:0] _T_2988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5597;
  reg [31:0] _T_2989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5598;
  reg [31:0] _T_2989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5599;
  reg [31:0] _T_2990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5600;
  reg [31:0] _T_2990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5601;
  reg [31:0] _T_2991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5602;
  reg [31:0] _T_2991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5603;
  reg [31:0] _T_2992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5604;
  reg [31:0] _T_2992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5605;
  reg [31:0] _T_2993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5606;
  reg [31:0] _T_2993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5607;
  reg [31:0] _T_2994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5608;
  reg [31:0] _T_2994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5609;
  reg [31:0] _T_2995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5610;
  reg [31:0] _T_2995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5611;
  reg [31:0] _T_2996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5612;
  reg [31:0] _T_2996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5613;
  reg [31:0] _T_2997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5614;
  reg [31:0] _T_2997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5615;
  reg [31:0] _T_2998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5616;
  reg [31:0] _T_2998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5617;
  reg [31:0] _T_2999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5618;
  reg [31:0] _T_2999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5619;
  reg [31:0] _T_3000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5620;
  reg [31:0] _T_3000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5621;
  reg [31:0] _T_3001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5622;
  reg [31:0] _T_3001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5623;
  reg [31:0] _T_3002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5624;
  reg [31:0] _T_3002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5625;
  reg [31:0] _T_3003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5626;
  reg [31:0] _T_3003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5627;
  reg [31:0] _T_3004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5628;
  reg [31:0] _T_3004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5629;
  reg [31:0] _T_3005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5630;
  reg [31:0] _T_3005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5631;
  reg [31:0] _T_3006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5632;
  reg [31:0] _T_3006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5633;
  reg [31:0] _T_3007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5634;
  reg [31:0] _T_3007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5635;
  reg [31:0] _T_3008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5636;
  reg [31:0] _T_3008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5637;
  reg [31:0] _T_3009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5638;
  reg [31:0] _T_3009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5639;
  reg [31:0] _T_3010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5640;
  reg [31:0] _T_3010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5641;
  reg [31:0] _T_3011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5642;
  reg [31:0] _T_3011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5643;
  reg [31:0] _T_3012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5644;
  reg [31:0] _T_3012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5645;
  reg [31:0] _T_3013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5646;
  reg [31:0] _T_3013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5647;
  reg [31:0] _T_3014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5648;
  reg [31:0] _T_3014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5649;
  reg [31:0] _T_3015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5650;
  reg [31:0] _T_3015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5651;
  reg [31:0] _T_3016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5652;
  reg [31:0] _T_3016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5653;
  reg [31:0] _T_3017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5654;
  reg [31:0] _T_3017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5655;
  reg [31:0] _T_3018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5656;
  reg [31:0] _T_3018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5657;
  reg [31:0] _T_3019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5658;
  reg [31:0] _T_3019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5659;
  reg [31:0] _T_3020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5660;
  reg [31:0] _T_3020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5661;
  reg [31:0] _T_3021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5662;
  reg [31:0] _T_3021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5663;
  reg [31:0] _T_3022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5664;
  reg [31:0] _T_3022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5665;
  reg [31:0] _T_3023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5666;
  reg [31:0] _T_3023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5667;
  reg [31:0] _T_3024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5668;
  reg [31:0] _T_3024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5669;
  reg [31:0] _T_3025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5670;
  reg [31:0] _T_3025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5671;
  reg [31:0] _T_3026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5672;
  reg [31:0] _T_3026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5673;
  reg [31:0] _T_3027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5674;
  reg [31:0] _T_3027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5675;
  reg [31:0] _T_3028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5676;
  reg [31:0] _T_3028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5677;
  reg [31:0] _T_3029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5678;
  reg [31:0] _T_3029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5679;
  reg [31:0] _T_3030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5680;
  reg [31:0] _T_3030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5681;
  reg [31:0] _T_3031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5682;
  reg [31:0] _T_3031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5683;
  reg [31:0] _T_3032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5684;
  reg [31:0] _T_3032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5685;
  reg [31:0] _T_3033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5686;
  reg [31:0] _T_3033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5687;
  reg [31:0] _T_3034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5688;
  reg [31:0] _T_3034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5689;
  reg [31:0] _T_3035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5690;
  reg [31:0] _T_3035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5691;
  reg [31:0] _T_3036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5692;
  reg [31:0] _T_3036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5693;
  reg [31:0] _T_3037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5694;
  reg [31:0] _T_3037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5695;
  reg [31:0] _T_3038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5696;
  reg [31:0] _T_3038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5697;
  reg [31:0] _T_3039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5698;
  reg [31:0] _T_3039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5699;
  reg [31:0] _T_3040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5700;
  reg [31:0] _T_3040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5701;
  reg [31:0] _T_3041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5702;
  reg [31:0] _T_3041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5703;
  reg [31:0] _T_3042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5704;
  reg [31:0] _T_3042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5705;
  reg [31:0] _T_3043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5706;
  reg [31:0] _T_3043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5707;
  reg [31:0] _T_3044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5708;
  reg [31:0] _T_3044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5709;
  reg [31:0] _T_3045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5710;
  reg [31:0] _T_3045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5711;
  reg [31:0] _T_3046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5712;
  reg [31:0] _T_3046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5713;
  reg [31:0] _T_3047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5714;
  reg [31:0] _T_3047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5715;
  reg [31:0] _T_3048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5716;
  reg [31:0] _T_3048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5717;
  reg [31:0] _T_3049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5718;
  reg [31:0] _T_3049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5719;
  reg [31:0] _T_3050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5720;
  reg [31:0] _T_3050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5721;
  reg [31:0] _T_3051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5722;
  reg [31:0] _T_3051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5723;
  reg [31:0] _T_3052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5724;
  reg [31:0] _T_3052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5725;
  reg [31:0] _T_3053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5726;
  reg [31:0] _T_3053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5727;
  reg [31:0] _T_3054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5728;
  reg [31:0] _T_3054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5729;
  reg [31:0] _T_3055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5730;
  reg [31:0] _T_3055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5731;
  reg [31:0] _T_3056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5732;
  reg [31:0] _T_3056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5733;
  reg [31:0] _T_3057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5734;
  reg [31:0] _T_3057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5735;
  reg [31:0] _T_3058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5736;
  reg [31:0] _T_3058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5737;
  reg [31:0] _T_3059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5738;
  reg [31:0] _T_3059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5739;
  reg [31:0] _T_3060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5740;
  reg [31:0] _T_3060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5741;
  reg [31:0] _T_3061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5742;
  reg [31:0] _T_3061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5743;
  reg [31:0] _T_3062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5744;
  reg [31:0] _T_3062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5745;
  reg [31:0] _T_3063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5746;
  reg [31:0] _T_3063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5747;
  reg [31:0] _T_3064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5748;
  reg [31:0] _T_3064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5749;
  reg [31:0] _T_3065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5750;
  reg [31:0] _T_3065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5751;
  reg [31:0] _T_3066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5752;
  reg [31:0] _T_3066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5753;
  reg [31:0] _T_3067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5754;
  reg [31:0] _T_3067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5755;
  reg [31:0] _T_3068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5756;
  reg [31:0] _T_3068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5757;
  reg [31:0] _T_3069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5758;
  reg [31:0] _T_3069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5759;
  reg [31:0] _T_3070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5760;
  reg [31:0] _T_3070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5761;
  reg [31:0] _T_3071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5762;
  reg [31:0] _T_3071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5763;
  reg [31:0] _T_3072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5764;
  reg [31:0] _T_3072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5765;
  reg [31:0] _T_3073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5766;
  reg [31:0] _T_3073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5767;
  reg [31:0] _T_3074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5768;
  reg [31:0] _T_3074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5769;
  reg [31:0] _T_3075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5770;
  reg [31:0] _T_3075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5771;
  reg [31:0] _T_3076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5772;
  reg [31:0] _T_3076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5773;
  reg [31:0] _T_3077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5774;
  reg [31:0] _T_3077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5775;
  reg [31:0] _T_3078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5776;
  reg [31:0] _T_3078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5777;
  reg [31:0] _T_3079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5778;
  reg [31:0] _T_3079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5779;
  reg [31:0] _T_3080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5780;
  reg [31:0] _T_3080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5781;
  reg [31:0] _T_3081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5782;
  reg [31:0] _T_3081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5783;
  reg [31:0] _T_3082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5784;
  reg [31:0] _T_3082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5785;
  reg [31:0] _T_3083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5786;
  reg [31:0] _T_3083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5787;
  reg [31:0] _T_3084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5788;
  reg [31:0] _T_3084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5789;
  reg [31:0] _T_3085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5790;
  reg [31:0] _T_3085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5791;
  reg [31:0] _T_3086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5792;
  reg [31:0] _T_3086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5793;
  reg [31:0] _T_3087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5794;
  reg [31:0] _T_3087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5795;
  reg [31:0] _T_3088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5796;
  reg [31:0] _T_3088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5797;
  reg [31:0] _T_3089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5798;
  reg [31:0] _T_3089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5799;
  reg [31:0] _T_3090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5800;
  reg [31:0] _T_3090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5801;
  reg [31:0] _T_3091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5802;
  reg [31:0] _T_3091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5803;
  reg [31:0] _T_3092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5804;
  reg [31:0] _T_3092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5805;
  reg [31:0] _T_3093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5806;
  reg [31:0] _T_3093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5807;
  reg [31:0] _T_3094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5808;
  reg [31:0] _T_3094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5809;
  reg [31:0] _T_3095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5810;
  reg [31:0] _T_3095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5811;
  reg [31:0] _T_3096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5812;
  reg [31:0] _T_3096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5813;
  reg [31:0] _T_3097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5814;
  reg [31:0] _T_3097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5815;
  reg [31:0] _T_3098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5816;
  reg [31:0] _T_3098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5817;
  reg [31:0] _T_3099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5818;
  reg [31:0] _T_3099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5819;
  reg [31:0] _T_3100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5820;
  reg [31:0] _T_3100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5821;
  reg [31:0] _T_3101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5822;
  reg [31:0] _T_3101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5823;
  reg [31:0] _T_3102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5824;
  reg [31:0] _T_3102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5825;
  reg [31:0] _T_3103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5826;
  reg [31:0] _T_3103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5827;
  reg [31:0] _T_3104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5828;
  reg [31:0] _T_3104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5829;
  reg [31:0] _T_3105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5830;
  reg [31:0] _T_3105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5831;
  reg [31:0] _T_3106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5832;
  reg [31:0] _T_3106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5833;
  reg [31:0] _T_3107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5834;
  reg [31:0] _T_3107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5835;
  reg [31:0] _T_3108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5836;
  reg [31:0] _T_3108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5837;
  reg [31:0] _T_3109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5838;
  reg [31:0] _T_3109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5839;
  reg [31:0] _T_3110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5840;
  reg [31:0] _T_3110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5841;
  reg [31:0] _T_3111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5842;
  reg [31:0] _T_3111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5843;
  reg [31:0] _T_3112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5844;
  reg [31:0] _T_3112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5845;
  reg [31:0] _T_3113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5846;
  reg [31:0] _T_3113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5847;
  reg [31:0] _T_3114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5848;
  reg [31:0] _T_3114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5849;
  reg [31:0] _T_3115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5850;
  reg [31:0] _T_3115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5851;
  reg [31:0] _T_3116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5852;
  reg [31:0] _T_3116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5853;
  reg [31:0] _T_3117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5854;
  reg [31:0] _T_3117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5855;
  reg [31:0] _T_3118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5856;
  reg [31:0] _T_3118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5857;
  reg [31:0] _T_3119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5858;
  reg [31:0] _T_3119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5859;
  reg [31:0] _T_3120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5860;
  reg [31:0] _T_3120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5861;
  reg [31:0] _T_3121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5862;
  reg [31:0] _T_3121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5863;
  reg [31:0] _T_3122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5864;
  reg [31:0] _T_3122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5865;
  reg [31:0] _T_3123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5866;
  reg [31:0] _T_3123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5867;
  reg [31:0] _T_3124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5868;
  reg [31:0] _T_3124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5869;
  reg [31:0] _T_3125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5870;
  reg [31:0] _T_3125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5871;
  reg [31:0] _T_3126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5872;
  reg [31:0] _T_3126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5873;
  reg [31:0] _T_3127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5874;
  reg [31:0] _T_3127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5875;
  reg [31:0] _T_3128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5876;
  reg [31:0] _T_3128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5877;
  reg [31:0] _T_3129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5878;
  reg [31:0] _T_3129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5879;
  reg [31:0] _T_3130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5880;
  reg [31:0] _T_3130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5881;
  reg [31:0] _T_3131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5882;
  reg [31:0] _T_3131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5883;
  reg [31:0] _T_3132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5884;
  reg [31:0] _T_3132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5885;
  reg [31:0] _T_3133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5886;
  reg [31:0] _T_3133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5887;
  reg [31:0] _T_3134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5888;
  reg [31:0] _T_3134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5889;
  reg [31:0] _T_3135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5890;
  reg [31:0] _T_3135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5891;
  reg [31:0] _T_3136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5892;
  reg [31:0] _T_3136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5893;
  reg [31:0] _T_3137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5894;
  reg [31:0] _T_3137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5895;
  reg [31:0] _T_3138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5896;
  reg [31:0] _T_3138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5897;
  reg [31:0] _T_3139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5898;
  reg [31:0] _T_3139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5899;
  reg [31:0] _T_3140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5900;
  reg [31:0] _T_3140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5901;
  reg [31:0] _T_3141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5902;
  reg [31:0] _T_3141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5903;
  reg [31:0] _T_3142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5904;
  reg [31:0] _T_3142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5905;
  reg [31:0] _T_3143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5906;
  reg [31:0] _T_3143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5907;
  reg [31:0] _T_3144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5908;
  reg [31:0] _T_3144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5909;
  reg [31:0] _T_3145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5910;
  reg [31:0] _T_3145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5911;
  reg [31:0] _T_3146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5912;
  reg [31:0] _T_3146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5913;
  reg [31:0] _T_3147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5914;
  reg [31:0] _T_3147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5915;
  reg [31:0] _T_3148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5916;
  reg [31:0] _T_3148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5917;
  reg [31:0] _T_3149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5918;
  reg [31:0] _T_3149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5919;
  reg [31:0] _T_3150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5920;
  reg [31:0] _T_3150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5921;
  reg [31:0] _T_3151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5922;
  reg [31:0] _T_3151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5923;
  reg [31:0] _T_3152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5924;
  reg [31:0] _T_3152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5925;
  reg [31:0] _T_3153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5926;
  reg [31:0] _T_3153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5927;
  reg [31:0] _T_3154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5928;
  reg [31:0] _T_3154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5929;
  reg [31:0] _T_3155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5930;
  reg [31:0] _T_3155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5931;
  reg [31:0] _T_3156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5932;
  reg [31:0] _T_3156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5933;
  reg [31:0] _T_3157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5934;
  reg [31:0] _T_3157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5935;
  reg [31:0] _T_3158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5936;
  reg [31:0] _T_3158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5937;
  reg [31:0] _T_3159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5938;
  reg [31:0] _T_3159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5939;
  reg [31:0] _T_3160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5940;
  reg [31:0] _T_3160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5941;
  reg [31:0] _T_3161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5942;
  reg [31:0] _T_3161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5943;
  reg [31:0] _T_3162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5944;
  reg [31:0] _T_3162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5945;
  reg [31:0] _T_3163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5946;
  reg [31:0] _T_3163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5947;
  reg [31:0] _T_3164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5948;
  reg [31:0] _T_3164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5949;
  reg [31:0] _T_3165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5950;
  reg [31:0] _T_3165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5951;
  reg [31:0] _T_3166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5952;
  reg [31:0] _T_3166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5953;
  reg [31:0] _T_3167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5954;
  reg [31:0] _T_3167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5955;
  reg [31:0] _T_3168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5956;
  reg [31:0] _T_3168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5957;
  reg [31:0] _T_3169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5958;
  reg [31:0] _T_3169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5959;
  reg [31:0] _T_3170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5960;
  reg [31:0] _T_3170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5961;
  reg [31:0] _T_3171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5962;
  reg [31:0] _T_3171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5963;
  reg [31:0] _T_3172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5964;
  reg [31:0] _T_3172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5965;
  reg [31:0] _T_3173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5966;
  reg [31:0] _T_3173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5967;
  reg [31:0] _T_3174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5968;
  reg [31:0] _T_3174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5969;
  reg [31:0] _T_3175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5970;
  reg [31:0] _T_3175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5971;
  reg [31:0] _T_3176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5972;
  reg [31:0] _T_3176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5973;
  reg [31:0] _T_3177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5974;
  reg [31:0] _T_3177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5975;
  reg [31:0] _T_3178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5976;
  reg [31:0] _T_3178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5977;
  reg [31:0] _T_3179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5978;
  reg [31:0] _T_3179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5979;
  reg [31:0] _T_3180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5980;
  reg [31:0] _T_3180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5981;
  reg [31:0] _T_3181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5982;
  reg [31:0] _T_3181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5983;
  reg [31:0] _T_3182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5984;
  reg [31:0] _T_3182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5985;
  reg [31:0] _T_3183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5986;
  reg [31:0] _T_3183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5987;
  reg [31:0] _T_3184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5988;
  reg [31:0] _T_3184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5989;
  reg [31:0] _T_3185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5990;
  reg [31:0] _T_3185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5991;
  reg [31:0] _T_3186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5992;
  reg [31:0] _T_3186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5993;
  reg [31:0] _T_3187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5994;
  reg [31:0] _T_3187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5995;
  reg [31:0] _T_3188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5996;
  reg [31:0] _T_3188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5997;
  reg [31:0] _T_3189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5998;
  reg [31:0] _T_3189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5999;
  reg [31:0] _T_3190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6000;
  reg [31:0] _T_3190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6001;
  reg [31:0] _T_3191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6002;
  reg [31:0] _T_3191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6003;
  reg [31:0] _T_3192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6004;
  reg [31:0] _T_3192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6005;
  reg [31:0] _T_3193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6006;
  reg [31:0] _T_3193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6007;
  reg [31:0] _T_3194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6008;
  reg [31:0] _T_3194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6009;
  reg [31:0] _T_3195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6010;
  reg [31:0] _T_3195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6011;
  reg [31:0] _T_3196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6012;
  reg [31:0] _T_3196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6013;
  reg [31:0] _T_3197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6014;
  reg [31:0] _T_3197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6015;
  reg [31:0] _T_3198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6016;
  reg [31:0] _T_3198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6017;
  reg [31:0] _T_3199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6018;
  reg [31:0] _T_3199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6019;
  reg [31:0] _T_3200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6020;
  reg [31:0] _T_3200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6021;
  reg [31:0] _T_3201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6022;
  reg [31:0] _T_3201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6023;
  reg [31:0] _T_3202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6024;
  reg [31:0] _T_3202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6025;
  reg [31:0] _T_3203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6026;
  reg [31:0] _T_3203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6027;
  reg [31:0] _T_3204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6028;
  reg [31:0] _T_3204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6029;
  reg [31:0] _T_3205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6030;
  reg [31:0] _T_3205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6031;
  reg [31:0] _T_3206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6032;
  reg [31:0] _T_3206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6033;
  reg [31:0] _T_3207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6034;
  reg [31:0] _T_3207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6035;
  reg [31:0] _T_3208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6036;
  reg [31:0] _T_3208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6037;
  reg [31:0] _T_3209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6038;
  reg [31:0] _T_3209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6039;
  reg [31:0] _T_3210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6040;
  reg [31:0] _T_3210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6041;
  reg [31:0] _T_3211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6042;
  reg [31:0] _T_3211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6043;
  reg [31:0] _T_3212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6044;
  reg [31:0] _T_3212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6045;
  reg [31:0] _T_3213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6046;
  reg [31:0] _T_3213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6047;
  reg [31:0] _T_3214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6048;
  reg [31:0] _T_3214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6049;
  reg [31:0] _T_3215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6050;
  reg [31:0] _T_3215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6051;
  reg [31:0] _T_3216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6052;
  reg [31:0] _T_3216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6053;
  reg [31:0] _T_3217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6054;
  reg [31:0] _T_3217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6055;
  reg [31:0] _T_3218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6056;
  reg [31:0] _T_3218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6057;
  reg [31:0] _T_3219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6058;
  reg [31:0] _T_3219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6059;
  reg [31:0] _T_3220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6060;
  reg [31:0] _T_3220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6061;
  reg [31:0] _T_3221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6062;
  reg [31:0] _T_3221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6063;
  reg [31:0] _T_3222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6064;
  reg [31:0] _T_3222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6065;
  reg [31:0] _T_3223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6066;
  reg [31:0] _T_3223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6067;
  reg [31:0] _T_3224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6068;
  reg [31:0] _T_3224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6069;
  reg [31:0] _T_3225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6070;
  reg [31:0] _T_3225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6071;
  reg [31:0] _T_3226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6072;
  reg [31:0] _T_3226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6073;
  reg [31:0] _T_3227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6074;
  reg [31:0] _T_3227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6075;
  reg [31:0] _T_3228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6076;
  reg [31:0] _T_3228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6077;
  reg [31:0] _T_3229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6078;
  reg [31:0] _T_3229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6079;
  reg [31:0] _T_3230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6080;
  reg [31:0] _T_3230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6081;
  reg [31:0] _T_3231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6082;
  reg [31:0] _T_3231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6083;
  reg [31:0] _T_3232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6084;
  reg [31:0] _T_3232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6085;
  reg [31:0] _T_3233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6086;
  reg [31:0] _T_3233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6087;
  reg [31:0] _T_3234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6088;
  reg [31:0] _T_3234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6089;
  reg [31:0] _T_3235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6090;
  reg [31:0] _T_3235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6091;
  reg [31:0] _T_3236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6092;
  reg [31:0] _T_3236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6093;
  reg [31:0] _T_3237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6094;
  reg [31:0] _T_3237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6095;
  reg [31:0] _T_3238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6096;
  reg [31:0] _T_3238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6097;
  reg [31:0] _T_3239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6098;
  reg [31:0] _T_3239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6099;
  reg [31:0] _T_3240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6100;
  reg [31:0] _T_3240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6101;
  reg [31:0] _T_3241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6102;
  reg [31:0] _T_3241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6103;
  reg [31:0] _T_3242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6104;
  reg [31:0] _T_3242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6105;
  reg [31:0] _T_3243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6106;
  reg [31:0] _T_3243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6107;
  reg [31:0] _T_3244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6108;
  reg [31:0] _T_3244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6109;
  reg [31:0] _T_3245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6110;
  reg [31:0] _T_3245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6111;
  reg [31:0] _T_3246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6112;
  reg [31:0] _T_3246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6113;
  reg [31:0] _T_3247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6114;
  reg [31:0] _T_3247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6115;
  reg [31:0] _T_3248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6116;
  reg [31:0] _T_3248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6117;
  reg [31:0] _T_3249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6118;
  reg [31:0] _T_3249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6119;
  reg [31:0] _T_3250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6120;
  reg [31:0] _T_3250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6121;
  reg [31:0] _T_3251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6122;
  reg [31:0] _T_3251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6123;
  reg [31:0] _T_3252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6124;
  reg [31:0] _T_3252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6125;
  reg [31:0] _T_3253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6126;
  reg [31:0] _T_3253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6127;
  reg [31:0] _T_3254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6128;
  reg [31:0] _T_3254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6129;
  reg [31:0] _T_3255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6130;
  reg [31:0] _T_3255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6131;
  reg [31:0] _T_3256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6132;
  reg [31:0] _T_3256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6133;
  reg [31:0] _T_3257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6134;
  reg [31:0] _T_3257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6135;
  reg [31:0] _T_3258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6136;
  reg [31:0] _T_3258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6137;
  reg [31:0] _T_3259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6138;
  reg [31:0] _T_3259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6139;
  reg [31:0] _T_3260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6140;
  reg [31:0] _T_3260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6141;
  reg [31:0] _T_3261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6142;
  reg [31:0] _T_3261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6143;
  reg [31:0] _T_3262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6144;
  reg [31:0] _T_3262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6145;
  wire [31:0] _GEN_10243 = 10'h2 == cnt[9:0] ? $signed(32'shffff) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10244 = 10'h3 == cnt[9:0] ? $signed(32'shfffd) : $signed(_GEN_10243); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10245 = 10'h4 == cnt[9:0] ? $signed(32'shfffb) : $signed(_GEN_10244); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10246 = 10'h5 == cnt[9:0] ? $signed(32'shfff8) : $signed(_GEN_10245); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10247 = 10'h6 == cnt[9:0] ? $signed(32'shfff5) : $signed(_GEN_10246); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10248 = 10'h7 == cnt[9:0] ? $signed(32'shfff1) : $signed(_GEN_10247); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10249 = 10'h8 == cnt[9:0] ? $signed(32'shffec) : $signed(_GEN_10248); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10250 = 10'h9 == cnt[9:0] ? $signed(32'shffe7) : $signed(_GEN_10249); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10251 = 10'ha == cnt[9:0] ? $signed(32'shffe1) : $signed(_GEN_10250); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10252 = 10'hb == cnt[9:0] ? $signed(32'shffdb) : $signed(_GEN_10251); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10253 = 10'hc == cnt[9:0] ? $signed(32'shffd4) : $signed(_GEN_10252); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10254 = 10'hd == cnt[9:0] ? $signed(32'shffcc) : $signed(_GEN_10253); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10255 = 10'he == cnt[9:0] ? $signed(32'shffc4) : $signed(_GEN_10254); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10256 = 10'hf == cnt[9:0] ? $signed(32'shffbb) : $signed(_GEN_10255); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10257 = 10'h10 == cnt[9:0] ? $signed(32'shffb1) : $signed(_GEN_10256); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10258 = 10'h11 == cnt[9:0] ? $signed(32'shffa7) : $signed(_GEN_10257); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10259 = 10'h12 == cnt[9:0] ? $signed(32'shff9c) : $signed(_GEN_10258); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10260 = 10'h13 == cnt[9:0] ? $signed(32'shff91) : $signed(_GEN_10259); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10261 = 10'h14 == cnt[9:0] ? $signed(32'shff85) : $signed(_GEN_10260); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10262 = 10'h15 == cnt[9:0] ? $signed(32'shff78) : $signed(_GEN_10261); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10263 = 10'h16 == cnt[9:0] ? $signed(32'shff6b) : $signed(_GEN_10262); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10264 = 10'h17 == cnt[9:0] ? $signed(32'shff5d) : $signed(_GEN_10263); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10265 = 10'h18 == cnt[9:0] ? $signed(32'shff4e) : $signed(_GEN_10264); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10266 = 10'h19 == cnt[9:0] ? $signed(32'shff3f) : $signed(_GEN_10265); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10267 = 10'h1a == cnt[9:0] ? $signed(32'shff30) : $signed(_GEN_10266); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10268 = 10'h1b == cnt[9:0] ? $signed(32'shff1f) : $signed(_GEN_10267); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10269 = 10'h1c == cnt[9:0] ? $signed(32'shff0e) : $signed(_GEN_10268); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10270 = 10'h1d == cnt[9:0] ? $signed(32'shfefd) : $signed(_GEN_10269); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10271 = 10'h1e == cnt[9:0] ? $signed(32'shfeeb) : $signed(_GEN_10270); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10272 = 10'h1f == cnt[9:0] ? $signed(32'shfed8) : $signed(_GEN_10271); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10273 = 10'h20 == cnt[9:0] ? $signed(32'shfec4) : $signed(_GEN_10272); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10274 = 10'h21 == cnt[9:0] ? $signed(32'shfeb0) : $signed(_GEN_10273); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10275 = 10'h22 == cnt[9:0] ? $signed(32'shfe9c) : $signed(_GEN_10274); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10276 = 10'h23 == cnt[9:0] ? $signed(32'shfe87) : $signed(_GEN_10275); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10277 = 10'h24 == cnt[9:0] ? $signed(32'shfe71) : $signed(_GEN_10276); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10278 = 10'h25 == cnt[9:0] ? $signed(32'shfe5a) : $signed(_GEN_10277); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10279 = 10'h26 == cnt[9:0] ? $signed(32'shfe43) : $signed(_GEN_10278); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10280 = 10'h27 == cnt[9:0] ? $signed(32'shfe2b) : $signed(_GEN_10279); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10281 = 10'h28 == cnt[9:0] ? $signed(32'shfe13) : $signed(_GEN_10280); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10282 = 10'h29 == cnt[9:0] ? $signed(32'shfdfa) : $signed(_GEN_10281); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10283 = 10'h2a == cnt[9:0] ? $signed(32'shfde1) : $signed(_GEN_10282); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10284 = 10'h2b == cnt[9:0] ? $signed(32'shfdc7) : $signed(_GEN_10283); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10285 = 10'h2c == cnt[9:0] ? $signed(32'shfdac) : $signed(_GEN_10284); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10286 = 10'h2d == cnt[9:0] ? $signed(32'shfd90) : $signed(_GEN_10285); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10287 = 10'h2e == cnt[9:0] ? $signed(32'shfd74) : $signed(_GEN_10286); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10288 = 10'h2f == cnt[9:0] ? $signed(32'shfd58) : $signed(_GEN_10287); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10289 = 10'h30 == cnt[9:0] ? $signed(32'shfd3b) : $signed(_GEN_10288); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10290 = 10'h31 == cnt[9:0] ? $signed(32'shfd1d) : $signed(_GEN_10289); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10291 = 10'h32 == cnt[9:0] ? $signed(32'shfcfe) : $signed(_GEN_10290); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10292 = 10'h33 == cnt[9:0] ? $signed(32'shfcdf) : $signed(_GEN_10291); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10293 = 10'h34 == cnt[9:0] ? $signed(32'shfcc0) : $signed(_GEN_10292); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10294 = 10'h35 == cnt[9:0] ? $signed(32'shfca0) : $signed(_GEN_10293); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10295 = 10'h36 == cnt[9:0] ? $signed(32'shfc7f) : $signed(_GEN_10294); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10296 = 10'h37 == cnt[9:0] ? $signed(32'shfc5d) : $signed(_GEN_10295); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10297 = 10'h38 == cnt[9:0] ? $signed(32'shfc3b) : $signed(_GEN_10296); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10298 = 10'h39 == cnt[9:0] ? $signed(32'shfc18) : $signed(_GEN_10297); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10299 = 10'h3a == cnt[9:0] ? $signed(32'shfbf5) : $signed(_GEN_10298); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10300 = 10'h3b == cnt[9:0] ? $signed(32'shfbd1) : $signed(_GEN_10299); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10301 = 10'h3c == cnt[9:0] ? $signed(32'shfbad) : $signed(_GEN_10300); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10302 = 10'h3d == cnt[9:0] ? $signed(32'shfb88) : $signed(_GEN_10301); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10303 = 10'h3e == cnt[9:0] ? $signed(32'shfb62) : $signed(_GEN_10302); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10304 = 10'h3f == cnt[9:0] ? $signed(32'shfb3c) : $signed(_GEN_10303); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10305 = 10'h40 == cnt[9:0] ? $signed(32'shfb15) : $signed(_GEN_10304); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10306 = 10'h41 == cnt[9:0] ? $signed(32'shfaed) : $signed(_GEN_10305); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10307 = 10'h42 == cnt[9:0] ? $signed(32'shfac5) : $signed(_GEN_10306); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10308 = 10'h43 == cnt[9:0] ? $signed(32'shfa9c) : $signed(_GEN_10307); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10309 = 10'h44 == cnt[9:0] ? $signed(32'shfa73) : $signed(_GEN_10308); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10310 = 10'h45 == cnt[9:0] ? $signed(32'shfa49) : $signed(_GEN_10309); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10311 = 10'h46 == cnt[9:0] ? $signed(32'shfa1f) : $signed(_GEN_10310); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10312 = 10'h47 == cnt[9:0] ? $signed(32'shf9f3) : $signed(_GEN_10311); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10313 = 10'h48 == cnt[9:0] ? $signed(32'shf9c8) : $signed(_GEN_10312); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10314 = 10'h49 == cnt[9:0] ? $signed(32'shf99b) : $signed(_GEN_10313); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10315 = 10'h4a == cnt[9:0] ? $signed(32'shf96e) : $signed(_GEN_10314); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10316 = 10'h4b == cnt[9:0] ? $signed(32'shf941) : $signed(_GEN_10315); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10317 = 10'h4c == cnt[9:0] ? $signed(32'shf913) : $signed(_GEN_10316); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10318 = 10'h4d == cnt[9:0] ? $signed(32'shf8e4) : $signed(_GEN_10317); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10319 = 10'h4e == cnt[9:0] ? $signed(32'shf8b4) : $signed(_GEN_10318); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10320 = 10'h4f == cnt[9:0] ? $signed(32'shf885) : $signed(_GEN_10319); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10321 = 10'h50 == cnt[9:0] ? $signed(32'shf854) : $signed(_GEN_10320); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10322 = 10'h51 == cnt[9:0] ? $signed(32'shf823) : $signed(_GEN_10321); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10323 = 10'h52 == cnt[9:0] ? $signed(32'shf7f1) : $signed(_GEN_10322); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10324 = 10'h53 == cnt[9:0] ? $signed(32'shf7bf) : $signed(_GEN_10323); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10325 = 10'h54 == cnt[9:0] ? $signed(32'shf78c) : $signed(_GEN_10324); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10326 = 10'h55 == cnt[9:0] ? $signed(32'shf758) : $signed(_GEN_10325); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10327 = 10'h56 == cnt[9:0] ? $signed(32'shf724) : $signed(_GEN_10326); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10328 = 10'h57 == cnt[9:0] ? $signed(32'shf6ef) : $signed(_GEN_10327); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10329 = 10'h58 == cnt[9:0] ? $signed(32'shf6ba) : $signed(_GEN_10328); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10330 = 10'h59 == cnt[9:0] ? $signed(32'shf684) : $signed(_GEN_10329); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10331 = 10'h5a == cnt[9:0] ? $signed(32'shf64e) : $signed(_GEN_10330); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10332 = 10'h5b == cnt[9:0] ? $signed(32'shf616) : $signed(_GEN_10331); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10333 = 10'h5c == cnt[9:0] ? $signed(32'shf5df) : $signed(_GEN_10332); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10334 = 10'h5d == cnt[9:0] ? $signed(32'shf5a6) : $signed(_GEN_10333); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10335 = 10'h5e == cnt[9:0] ? $signed(32'shf56e) : $signed(_GEN_10334); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10336 = 10'h5f == cnt[9:0] ? $signed(32'shf534) : $signed(_GEN_10335); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10337 = 10'h60 == cnt[9:0] ? $signed(32'shf4fa) : $signed(_GEN_10336); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10338 = 10'h61 == cnt[9:0] ? $signed(32'shf4bf) : $signed(_GEN_10337); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10339 = 10'h62 == cnt[9:0] ? $signed(32'shf484) : $signed(_GEN_10338); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10340 = 10'h63 == cnt[9:0] ? $signed(32'shf448) : $signed(_GEN_10339); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10341 = 10'h64 == cnt[9:0] ? $signed(32'shf40c) : $signed(_GEN_10340); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10342 = 10'h65 == cnt[9:0] ? $signed(32'shf3cf) : $signed(_GEN_10341); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10343 = 10'h66 == cnt[9:0] ? $signed(32'shf391) : $signed(_GEN_10342); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10344 = 10'h67 == cnt[9:0] ? $signed(32'shf353) : $signed(_GEN_10343); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10345 = 10'h68 == cnt[9:0] ? $signed(32'shf314) : $signed(_GEN_10344); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10346 = 10'h69 == cnt[9:0] ? $signed(32'shf2d5) : $signed(_GEN_10345); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10347 = 10'h6a == cnt[9:0] ? $signed(32'shf295) : $signed(_GEN_10346); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10348 = 10'h6b == cnt[9:0] ? $signed(32'shf254) : $signed(_GEN_10347); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10349 = 10'h6c == cnt[9:0] ? $signed(32'shf213) : $signed(_GEN_10348); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10350 = 10'h6d == cnt[9:0] ? $signed(32'shf1d2) : $signed(_GEN_10349); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10351 = 10'h6e == cnt[9:0] ? $signed(32'shf18f) : $signed(_GEN_10350); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10352 = 10'h6f == cnt[9:0] ? $signed(32'shf14c) : $signed(_GEN_10351); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10353 = 10'h70 == cnt[9:0] ? $signed(32'shf109) : $signed(_GEN_10352); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10354 = 10'h71 == cnt[9:0] ? $signed(32'shf0c5) : $signed(_GEN_10353); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10355 = 10'h72 == cnt[9:0] ? $signed(32'shf080) : $signed(_GEN_10354); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10356 = 10'h73 == cnt[9:0] ? $signed(32'shf03b) : $signed(_GEN_10355); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10357 = 10'h74 == cnt[9:0] ? $signed(32'sheff5) : $signed(_GEN_10356); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10358 = 10'h75 == cnt[9:0] ? $signed(32'shefaf) : $signed(_GEN_10357); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10359 = 10'h76 == cnt[9:0] ? $signed(32'shef68) : $signed(_GEN_10358); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10360 = 10'h77 == cnt[9:0] ? $signed(32'shef21) : $signed(_GEN_10359); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10361 = 10'h78 == cnt[9:0] ? $signed(32'sheed9) : $signed(_GEN_10360); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10362 = 10'h79 == cnt[9:0] ? $signed(32'shee90) : $signed(_GEN_10361); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10363 = 10'h7a == cnt[9:0] ? $signed(32'shee47) : $signed(_GEN_10362); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10364 = 10'h7b == cnt[9:0] ? $signed(32'shedfd) : $signed(_GEN_10363); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10365 = 10'h7c == cnt[9:0] ? $signed(32'shedb3) : $signed(_GEN_10364); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10366 = 10'h7d == cnt[9:0] ? $signed(32'shed68) : $signed(_GEN_10365); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10367 = 10'h7e == cnt[9:0] ? $signed(32'shed1c) : $signed(_GEN_10366); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10368 = 10'h7f == cnt[9:0] ? $signed(32'shecd0) : $signed(_GEN_10367); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10369 = 10'h80 == cnt[9:0] ? $signed(32'shec83) : $signed(_GEN_10368); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10370 = 10'h81 == cnt[9:0] ? $signed(32'shec36) : $signed(_GEN_10369); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10371 = 10'h82 == cnt[9:0] ? $signed(32'shebe8) : $signed(_GEN_10370); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10372 = 10'h83 == cnt[9:0] ? $signed(32'sheb9a) : $signed(_GEN_10371); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10373 = 10'h84 == cnt[9:0] ? $signed(32'sheb4b) : $signed(_GEN_10372); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10374 = 10'h85 == cnt[9:0] ? $signed(32'sheafc) : $signed(_GEN_10373); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10375 = 10'h86 == cnt[9:0] ? $signed(32'sheaab) : $signed(_GEN_10374); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10376 = 10'h87 == cnt[9:0] ? $signed(32'shea5b) : $signed(_GEN_10375); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10377 = 10'h88 == cnt[9:0] ? $signed(32'shea0a) : $signed(_GEN_10376); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10378 = 10'h89 == cnt[9:0] ? $signed(32'she9b8) : $signed(_GEN_10377); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10379 = 10'h8a == cnt[9:0] ? $signed(32'she966) : $signed(_GEN_10378); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10380 = 10'h8b == cnt[9:0] ? $signed(32'she913) : $signed(_GEN_10379); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10381 = 10'h8c == cnt[9:0] ? $signed(32'she8bf) : $signed(_GEN_10380); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10382 = 10'h8d == cnt[9:0] ? $signed(32'she86b) : $signed(_GEN_10381); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10383 = 10'h8e == cnt[9:0] ? $signed(32'she817) : $signed(_GEN_10382); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10384 = 10'h8f == cnt[9:0] ? $signed(32'she7c2) : $signed(_GEN_10383); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10385 = 10'h90 == cnt[9:0] ? $signed(32'she76c) : $signed(_GEN_10384); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10386 = 10'h91 == cnt[9:0] ? $signed(32'she716) : $signed(_GEN_10385); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10387 = 10'h92 == cnt[9:0] ? $signed(32'she6bf) : $signed(_GEN_10386); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10388 = 10'h93 == cnt[9:0] ? $signed(32'she667) : $signed(_GEN_10387); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10389 = 10'h94 == cnt[9:0] ? $signed(32'she610) : $signed(_GEN_10388); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10390 = 10'h95 == cnt[9:0] ? $signed(32'she5b7) : $signed(_GEN_10389); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10391 = 10'h96 == cnt[9:0] ? $signed(32'she55e) : $signed(_GEN_10390); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10392 = 10'h97 == cnt[9:0] ? $signed(32'she504) : $signed(_GEN_10391); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10393 = 10'h98 == cnt[9:0] ? $signed(32'she4aa) : $signed(_GEN_10392); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10394 = 10'h99 == cnt[9:0] ? $signed(32'she450) : $signed(_GEN_10393); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10395 = 10'h9a == cnt[9:0] ? $signed(32'she3f4) : $signed(_GEN_10394); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10396 = 10'h9b == cnt[9:0] ? $signed(32'she399) : $signed(_GEN_10395); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10397 = 10'h9c == cnt[9:0] ? $signed(32'she33c) : $signed(_GEN_10396); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10398 = 10'h9d == cnt[9:0] ? $signed(32'she2df) : $signed(_GEN_10397); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10399 = 10'h9e == cnt[9:0] ? $signed(32'she282) : $signed(_GEN_10398); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10400 = 10'h9f == cnt[9:0] ? $signed(32'she224) : $signed(_GEN_10399); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10401 = 10'ha0 == cnt[9:0] ? $signed(32'she1c6) : $signed(_GEN_10400); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10402 = 10'ha1 == cnt[9:0] ? $signed(32'she167) : $signed(_GEN_10401); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10403 = 10'ha2 == cnt[9:0] ? $signed(32'she107) : $signed(_GEN_10402); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10404 = 10'ha3 == cnt[9:0] ? $signed(32'she0a7) : $signed(_GEN_10403); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10405 = 10'ha4 == cnt[9:0] ? $signed(32'she046) : $signed(_GEN_10404); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10406 = 10'ha5 == cnt[9:0] ? $signed(32'shdfe5) : $signed(_GEN_10405); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10407 = 10'ha6 == cnt[9:0] ? $signed(32'shdf83) : $signed(_GEN_10406); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10408 = 10'ha7 == cnt[9:0] ? $signed(32'shdf21) : $signed(_GEN_10407); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10409 = 10'ha8 == cnt[9:0] ? $signed(32'shdebe) : $signed(_GEN_10408); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10410 = 10'ha9 == cnt[9:0] ? $signed(32'shde5b) : $signed(_GEN_10409); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10411 = 10'haa == cnt[9:0] ? $signed(32'shddf7) : $signed(_GEN_10410); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10412 = 10'hab == cnt[9:0] ? $signed(32'shdd92) : $signed(_GEN_10411); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10413 = 10'hac == cnt[9:0] ? $signed(32'shdd2d) : $signed(_GEN_10412); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10414 = 10'had == cnt[9:0] ? $signed(32'shdcc8) : $signed(_GEN_10413); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10415 = 10'hae == cnt[9:0] ? $signed(32'shdc62) : $signed(_GEN_10414); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10416 = 10'haf == cnt[9:0] ? $signed(32'shdbfb) : $signed(_GEN_10415); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10417 = 10'hb0 == cnt[9:0] ? $signed(32'shdb94) : $signed(_GEN_10416); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10418 = 10'hb1 == cnt[9:0] ? $signed(32'shdb2c) : $signed(_GEN_10417); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10419 = 10'hb2 == cnt[9:0] ? $signed(32'shdac4) : $signed(_GEN_10418); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10420 = 10'hb3 == cnt[9:0] ? $signed(32'shda5c) : $signed(_GEN_10419); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10421 = 10'hb4 == cnt[9:0] ? $signed(32'shd9f2) : $signed(_GEN_10420); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10422 = 10'hb5 == cnt[9:0] ? $signed(32'shd989) : $signed(_GEN_10421); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10423 = 10'hb6 == cnt[9:0] ? $signed(32'shd91e) : $signed(_GEN_10422); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10424 = 10'hb7 == cnt[9:0] ? $signed(32'shd8b4) : $signed(_GEN_10423); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10425 = 10'hb8 == cnt[9:0] ? $signed(32'shd848) : $signed(_GEN_10424); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10426 = 10'hb9 == cnt[9:0] ? $signed(32'shd7dc) : $signed(_GEN_10425); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10427 = 10'hba == cnt[9:0] ? $signed(32'shd770) : $signed(_GEN_10426); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10428 = 10'hbb == cnt[9:0] ? $signed(32'shd703) : $signed(_GEN_10427); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10429 = 10'hbc == cnt[9:0] ? $signed(32'shd696) : $signed(_GEN_10428); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10430 = 10'hbd == cnt[9:0] ? $signed(32'shd628) : $signed(_GEN_10429); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10431 = 10'hbe == cnt[9:0] ? $signed(32'shd5ba) : $signed(_GEN_10430); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10432 = 10'hbf == cnt[9:0] ? $signed(32'shd54b) : $signed(_GEN_10431); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10433 = 10'hc0 == cnt[9:0] ? $signed(32'shd4db) : $signed(_GEN_10432); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10434 = 10'hc1 == cnt[9:0] ? $signed(32'shd46b) : $signed(_GEN_10433); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10435 = 10'hc2 == cnt[9:0] ? $signed(32'shd3fb) : $signed(_GEN_10434); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10436 = 10'hc3 == cnt[9:0] ? $signed(32'shd38a) : $signed(_GEN_10435); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10437 = 10'hc4 == cnt[9:0] ? $signed(32'shd318) : $signed(_GEN_10436); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10438 = 10'hc5 == cnt[9:0] ? $signed(32'shd2a6) : $signed(_GEN_10437); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10439 = 10'hc6 == cnt[9:0] ? $signed(32'shd234) : $signed(_GEN_10438); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10440 = 10'hc7 == cnt[9:0] ? $signed(32'shd1c1) : $signed(_GEN_10439); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10441 = 10'hc8 == cnt[9:0] ? $signed(32'shd14d) : $signed(_GEN_10440); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10442 = 10'hc9 == cnt[9:0] ? $signed(32'shd0d9) : $signed(_GEN_10441); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10443 = 10'hca == cnt[9:0] ? $signed(32'shd065) : $signed(_GEN_10442); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10444 = 10'hcb == cnt[9:0] ? $signed(32'shcff0) : $signed(_GEN_10443); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10445 = 10'hcc == cnt[9:0] ? $signed(32'shcf7a) : $signed(_GEN_10444); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10446 = 10'hcd == cnt[9:0] ? $signed(32'shcf04) : $signed(_GEN_10445); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10447 = 10'hce == cnt[9:0] ? $signed(32'shce8e) : $signed(_GEN_10446); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10448 = 10'hcf == cnt[9:0] ? $signed(32'shce17) : $signed(_GEN_10447); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10449 = 10'hd0 == cnt[9:0] ? $signed(32'shcd9f) : $signed(_GEN_10448); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10450 = 10'hd1 == cnt[9:0] ? $signed(32'shcd27) : $signed(_GEN_10449); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10451 = 10'hd2 == cnt[9:0] ? $signed(32'shccae) : $signed(_GEN_10450); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10452 = 10'hd3 == cnt[9:0] ? $signed(32'shcc35) : $signed(_GEN_10451); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10453 = 10'hd4 == cnt[9:0] ? $signed(32'shcbbc) : $signed(_GEN_10452); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10454 = 10'hd5 == cnt[9:0] ? $signed(32'shcb42) : $signed(_GEN_10453); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10455 = 10'hd6 == cnt[9:0] ? $signed(32'shcac7) : $signed(_GEN_10454); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10456 = 10'hd7 == cnt[9:0] ? $signed(32'shca4d) : $signed(_GEN_10455); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10457 = 10'hd8 == cnt[9:0] ? $signed(32'shc9d1) : $signed(_GEN_10456); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10458 = 10'hd9 == cnt[9:0] ? $signed(32'shc955) : $signed(_GEN_10457); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10459 = 10'hda == cnt[9:0] ? $signed(32'shc8d9) : $signed(_GEN_10458); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10460 = 10'hdb == cnt[9:0] ? $signed(32'shc85c) : $signed(_GEN_10459); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10461 = 10'hdc == cnt[9:0] ? $signed(32'shc7de) : $signed(_GEN_10460); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10462 = 10'hdd == cnt[9:0] ? $signed(32'shc761) : $signed(_GEN_10461); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10463 = 10'hde == cnt[9:0] ? $signed(32'shc6e2) : $signed(_GEN_10462); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10464 = 10'hdf == cnt[9:0] ? $signed(32'shc663) : $signed(_GEN_10463); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10465 = 10'he0 == cnt[9:0] ? $signed(32'shc5e4) : $signed(_GEN_10464); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10466 = 10'he1 == cnt[9:0] ? $signed(32'shc564) : $signed(_GEN_10465); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10467 = 10'he2 == cnt[9:0] ? $signed(32'shc4e4) : $signed(_GEN_10466); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10468 = 10'he3 == cnt[9:0] ? $signed(32'shc463) : $signed(_GEN_10467); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10469 = 10'he4 == cnt[9:0] ? $signed(32'shc3e2) : $signed(_GEN_10468); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10470 = 10'he5 == cnt[9:0] ? $signed(32'shc360) : $signed(_GEN_10469); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10471 = 10'he6 == cnt[9:0] ? $signed(32'shc2de) : $signed(_GEN_10470); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10472 = 10'he7 == cnt[9:0] ? $signed(32'shc25c) : $signed(_GEN_10471); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10473 = 10'he8 == cnt[9:0] ? $signed(32'shc1d8) : $signed(_GEN_10472); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10474 = 10'he9 == cnt[9:0] ? $signed(32'shc155) : $signed(_GEN_10473); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10475 = 10'hea == cnt[9:0] ? $signed(32'shc0d1) : $signed(_GEN_10474); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10476 = 10'heb == cnt[9:0] ? $signed(32'shc04c) : $signed(_GEN_10475); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10477 = 10'hec == cnt[9:0] ? $signed(32'shbfc7) : $signed(_GEN_10476); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10478 = 10'hed == cnt[9:0] ? $signed(32'shbf42) : $signed(_GEN_10477); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10479 = 10'hee == cnt[9:0] ? $signed(32'shbebc) : $signed(_GEN_10478); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10480 = 10'hef == cnt[9:0] ? $signed(32'shbe36) : $signed(_GEN_10479); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10481 = 10'hf0 == cnt[9:0] ? $signed(32'shbdaf) : $signed(_GEN_10480); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10482 = 10'hf1 == cnt[9:0] ? $signed(32'shbd28) : $signed(_GEN_10481); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10483 = 10'hf2 == cnt[9:0] ? $signed(32'shbca0) : $signed(_GEN_10482); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10484 = 10'hf3 == cnt[9:0] ? $signed(32'shbc18) : $signed(_GEN_10483); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10485 = 10'hf4 == cnt[9:0] ? $signed(32'shbb8f) : $signed(_GEN_10484); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10486 = 10'hf5 == cnt[9:0] ? $signed(32'shbb06) : $signed(_GEN_10485); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10487 = 10'hf6 == cnt[9:0] ? $signed(32'shba7d) : $signed(_GEN_10486); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10488 = 10'hf7 == cnt[9:0] ? $signed(32'shb9f3) : $signed(_GEN_10487); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10489 = 10'hf8 == cnt[9:0] ? $signed(32'shb968) : $signed(_GEN_10488); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10490 = 10'hf9 == cnt[9:0] ? $signed(32'shb8dd) : $signed(_GEN_10489); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10491 = 10'hfa == cnt[9:0] ? $signed(32'shb852) : $signed(_GEN_10490); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10492 = 10'hfb == cnt[9:0] ? $signed(32'shb7c6) : $signed(_GEN_10491); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10493 = 10'hfc == cnt[9:0] ? $signed(32'shb73a) : $signed(_GEN_10492); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10494 = 10'hfd == cnt[9:0] ? $signed(32'shb6ad) : $signed(_GEN_10493); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10495 = 10'hfe == cnt[9:0] ? $signed(32'shb620) : $signed(_GEN_10494); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10496 = 10'hff == cnt[9:0] ? $signed(32'shb593) : $signed(_GEN_10495); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10497 = 10'h100 == cnt[9:0] ? $signed(32'shb505) : $signed(_GEN_10496); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10498 = 10'h101 == cnt[9:0] ? $signed(32'shb477) : $signed(_GEN_10497); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10499 = 10'h102 == cnt[9:0] ? $signed(32'shb3e8) : $signed(_GEN_10498); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10500 = 10'h103 == cnt[9:0] ? $signed(32'shb358) : $signed(_GEN_10499); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10501 = 10'h104 == cnt[9:0] ? $signed(32'shb2c9) : $signed(_GEN_10500); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10502 = 10'h105 == cnt[9:0] ? $signed(32'shb239) : $signed(_GEN_10501); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10503 = 10'h106 == cnt[9:0] ? $signed(32'shb1a8) : $signed(_GEN_10502); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10504 = 10'h107 == cnt[9:0] ? $signed(32'shb117) : $signed(_GEN_10503); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10505 = 10'h108 == cnt[9:0] ? $signed(32'shb086) : $signed(_GEN_10504); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10506 = 10'h109 == cnt[9:0] ? $signed(32'shaff4) : $signed(_GEN_10505); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10507 = 10'h10a == cnt[9:0] ? $signed(32'shaf62) : $signed(_GEN_10506); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10508 = 10'h10b == cnt[9:0] ? $signed(32'shaecf) : $signed(_GEN_10507); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10509 = 10'h10c == cnt[9:0] ? $signed(32'shae3c) : $signed(_GEN_10508); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10510 = 10'h10d == cnt[9:0] ? $signed(32'shada8) : $signed(_GEN_10509); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10511 = 10'h10e == cnt[9:0] ? $signed(32'shad14) : $signed(_GEN_10510); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10512 = 10'h10f == cnt[9:0] ? $signed(32'shac80) : $signed(_GEN_10511); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10513 = 10'h110 == cnt[9:0] ? $signed(32'shabeb) : $signed(_GEN_10512); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10514 = 10'h111 == cnt[9:0] ? $signed(32'shab56) : $signed(_GEN_10513); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10515 = 10'h112 == cnt[9:0] ? $signed(32'shaac1) : $signed(_GEN_10514); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10516 = 10'h113 == cnt[9:0] ? $signed(32'shaa2a) : $signed(_GEN_10515); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10517 = 10'h114 == cnt[9:0] ? $signed(32'sha994) : $signed(_GEN_10516); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10518 = 10'h115 == cnt[9:0] ? $signed(32'sha8fd) : $signed(_GEN_10517); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10519 = 10'h116 == cnt[9:0] ? $signed(32'sha866) : $signed(_GEN_10518); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10520 = 10'h117 == cnt[9:0] ? $signed(32'sha7ce) : $signed(_GEN_10519); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10521 = 10'h118 == cnt[9:0] ? $signed(32'sha736) : $signed(_GEN_10520); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10522 = 10'h119 == cnt[9:0] ? $signed(32'sha69e) : $signed(_GEN_10521); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10523 = 10'h11a == cnt[9:0] ? $signed(32'sha605) : $signed(_GEN_10522); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10524 = 10'h11b == cnt[9:0] ? $signed(32'sha56c) : $signed(_GEN_10523); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10525 = 10'h11c == cnt[9:0] ? $signed(32'sha4d2) : $signed(_GEN_10524); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10526 = 10'h11d == cnt[9:0] ? $signed(32'sha438) : $signed(_GEN_10525); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10527 = 10'h11e == cnt[9:0] ? $signed(32'sha39e) : $signed(_GEN_10526); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10528 = 10'h11f == cnt[9:0] ? $signed(32'sha303) : $signed(_GEN_10527); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10529 = 10'h120 == cnt[9:0] ? $signed(32'sha268) : $signed(_GEN_10528); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10530 = 10'h121 == cnt[9:0] ? $signed(32'sha1cc) : $signed(_GEN_10529); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10531 = 10'h122 == cnt[9:0] ? $signed(32'sha130) : $signed(_GEN_10530); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10532 = 10'h123 == cnt[9:0] ? $signed(32'sha094) : $signed(_GEN_10531); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10533 = 10'h124 == cnt[9:0] ? $signed(32'sh9ff7) : $signed(_GEN_10532); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10534 = 10'h125 == cnt[9:0] ? $signed(32'sh9f5a) : $signed(_GEN_10533); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10535 = 10'h126 == cnt[9:0] ? $signed(32'sh9ebc) : $signed(_GEN_10534); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10536 = 10'h127 == cnt[9:0] ? $signed(32'sh9e1e) : $signed(_GEN_10535); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10537 = 10'h128 == cnt[9:0] ? $signed(32'sh9d80) : $signed(_GEN_10536); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10538 = 10'h129 == cnt[9:0] ? $signed(32'sh9ce1) : $signed(_GEN_10537); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10539 = 10'h12a == cnt[9:0] ? $signed(32'sh9c42) : $signed(_GEN_10538); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10540 = 10'h12b == cnt[9:0] ? $signed(32'sh9ba3) : $signed(_GEN_10539); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10541 = 10'h12c == cnt[9:0] ? $signed(32'sh9b03) : $signed(_GEN_10540); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10542 = 10'h12d == cnt[9:0] ? $signed(32'sh9a63) : $signed(_GEN_10541); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10543 = 10'h12e == cnt[9:0] ? $signed(32'sh99c2) : $signed(_GEN_10542); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10544 = 10'h12f == cnt[9:0] ? $signed(32'sh9921) : $signed(_GEN_10543); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10545 = 10'h130 == cnt[9:0] ? $signed(32'sh9880) : $signed(_GEN_10544); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10546 = 10'h131 == cnt[9:0] ? $signed(32'sh97de) : $signed(_GEN_10545); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10547 = 10'h132 == cnt[9:0] ? $signed(32'sh973c) : $signed(_GEN_10546); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10548 = 10'h133 == cnt[9:0] ? $signed(32'sh969a) : $signed(_GEN_10547); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10549 = 10'h134 == cnt[9:0] ? $signed(32'sh95f7) : $signed(_GEN_10548); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10550 = 10'h135 == cnt[9:0] ? $signed(32'sh9554) : $signed(_GEN_10549); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10551 = 10'h136 == cnt[9:0] ? $signed(32'sh94b0) : $signed(_GEN_10550); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10552 = 10'h137 == cnt[9:0] ? $signed(32'sh940c) : $signed(_GEN_10551); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10553 = 10'h138 == cnt[9:0] ? $signed(32'sh9368) : $signed(_GEN_10552); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10554 = 10'h139 == cnt[9:0] ? $signed(32'sh92c4) : $signed(_GEN_10553); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10555 = 10'h13a == cnt[9:0] ? $signed(32'sh921f) : $signed(_GEN_10554); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10556 = 10'h13b == cnt[9:0] ? $signed(32'sh9179) : $signed(_GEN_10555); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10557 = 10'h13c == cnt[9:0] ? $signed(32'sh90d4) : $signed(_GEN_10556); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10558 = 10'h13d == cnt[9:0] ? $signed(32'sh902e) : $signed(_GEN_10557); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10559 = 10'h13e == cnt[9:0] ? $signed(32'sh8f88) : $signed(_GEN_10558); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10560 = 10'h13f == cnt[9:0] ? $signed(32'sh8ee1) : $signed(_GEN_10559); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10561 = 10'h140 == cnt[9:0] ? $signed(32'sh8e3a) : $signed(_GEN_10560); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10562 = 10'h141 == cnt[9:0] ? $signed(32'sh8d93) : $signed(_GEN_10561); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10563 = 10'h142 == cnt[9:0] ? $signed(32'sh8ceb) : $signed(_GEN_10562); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10564 = 10'h143 == cnt[9:0] ? $signed(32'sh8c43) : $signed(_GEN_10563); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10565 = 10'h144 == cnt[9:0] ? $signed(32'sh8b9a) : $signed(_GEN_10564); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10566 = 10'h145 == cnt[9:0] ? $signed(32'sh8af2) : $signed(_GEN_10565); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10567 = 10'h146 == cnt[9:0] ? $signed(32'sh8a49) : $signed(_GEN_10566); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10568 = 10'h147 == cnt[9:0] ? $signed(32'sh899f) : $signed(_GEN_10567); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10569 = 10'h148 == cnt[9:0] ? $signed(32'sh88f6) : $signed(_GEN_10568); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10570 = 10'h149 == cnt[9:0] ? $signed(32'sh884c) : $signed(_GEN_10569); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10571 = 10'h14a == cnt[9:0] ? $signed(32'sh87a1) : $signed(_GEN_10570); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10572 = 10'h14b == cnt[9:0] ? $signed(32'sh86f7) : $signed(_GEN_10571); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10573 = 10'h14c == cnt[9:0] ? $signed(32'sh864c) : $signed(_GEN_10572); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10574 = 10'h14d == cnt[9:0] ? $signed(32'sh85a0) : $signed(_GEN_10573); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10575 = 10'h14e == cnt[9:0] ? $signed(32'sh84f5) : $signed(_GEN_10574); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10576 = 10'h14f == cnt[9:0] ? $signed(32'sh8449) : $signed(_GEN_10575); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10577 = 10'h150 == cnt[9:0] ? $signed(32'sh839c) : $signed(_GEN_10576); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10578 = 10'h151 == cnt[9:0] ? $signed(32'sh82f0) : $signed(_GEN_10577); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10579 = 10'h152 == cnt[9:0] ? $signed(32'sh8243) : $signed(_GEN_10578); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10580 = 10'h153 == cnt[9:0] ? $signed(32'sh8195) : $signed(_GEN_10579); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10581 = 10'h154 == cnt[9:0] ? $signed(32'sh80e8) : $signed(_GEN_10580); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10582 = 10'h155 == cnt[9:0] ? $signed(32'sh803a) : $signed(_GEN_10581); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10583 = 10'h156 == cnt[9:0] ? $signed(32'sh7f8c) : $signed(_GEN_10582); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10584 = 10'h157 == cnt[9:0] ? $signed(32'sh7edd) : $signed(_GEN_10583); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10585 = 10'h158 == cnt[9:0] ? $signed(32'sh7e2f) : $signed(_GEN_10584); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10586 = 10'h159 == cnt[9:0] ? $signed(32'sh7d7f) : $signed(_GEN_10585); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10587 = 10'h15a == cnt[9:0] ? $signed(32'sh7cd0) : $signed(_GEN_10586); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10588 = 10'h15b == cnt[9:0] ? $signed(32'sh7c20) : $signed(_GEN_10587); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10589 = 10'h15c == cnt[9:0] ? $signed(32'sh7b70) : $signed(_GEN_10588); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10590 = 10'h15d == cnt[9:0] ? $signed(32'sh7ac0) : $signed(_GEN_10589); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10591 = 10'h15e == cnt[9:0] ? $signed(32'sh7a10) : $signed(_GEN_10590); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10592 = 10'h15f == cnt[9:0] ? $signed(32'sh795f) : $signed(_GEN_10591); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10593 = 10'h160 == cnt[9:0] ? $signed(32'sh78ad) : $signed(_GEN_10592); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10594 = 10'h161 == cnt[9:0] ? $signed(32'sh77fc) : $signed(_GEN_10593); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10595 = 10'h162 == cnt[9:0] ? $signed(32'sh774a) : $signed(_GEN_10594); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10596 = 10'h163 == cnt[9:0] ? $signed(32'sh7698) : $signed(_GEN_10595); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10597 = 10'h164 == cnt[9:0] ? $signed(32'sh75e6) : $signed(_GEN_10596); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10598 = 10'h165 == cnt[9:0] ? $signed(32'sh7533) : $signed(_GEN_10597); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10599 = 10'h166 == cnt[9:0] ? $signed(32'sh7480) : $signed(_GEN_10598); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10600 = 10'h167 == cnt[9:0] ? $signed(32'sh73cd) : $signed(_GEN_10599); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10601 = 10'h168 == cnt[9:0] ? $signed(32'sh731a) : $signed(_GEN_10600); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10602 = 10'h169 == cnt[9:0] ? $signed(32'sh7266) : $signed(_GEN_10601); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10603 = 10'h16a == cnt[9:0] ? $signed(32'sh71b2) : $signed(_GEN_10602); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10604 = 10'h16b == cnt[9:0] ? $signed(32'sh70fe) : $signed(_GEN_10603); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10605 = 10'h16c == cnt[9:0] ? $signed(32'sh7049) : $signed(_GEN_10604); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10606 = 10'h16d == cnt[9:0] ? $signed(32'sh6f94) : $signed(_GEN_10605); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10607 = 10'h16e == cnt[9:0] ? $signed(32'sh6edf) : $signed(_GEN_10606); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10608 = 10'h16f == cnt[9:0] ? $signed(32'sh6e2a) : $signed(_GEN_10607); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10609 = 10'h170 == cnt[9:0] ? $signed(32'sh6d74) : $signed(_GEN_10608); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10610 = 10'h171 == cnt[9:0] ? $signed(32'sh6cbe) : $signed(_GEN_10609); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10611 = 10'h172 == cnt[9:0] ? $signed(32'sh6c08) : $signed(_GEN_10610); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10612 = 10'h173 == cnt[9:0] ? $signed(32'sh6b52) : $signed(_GEN_10611); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10613 = 10'h174 == cnt[9:0] ? $signed(32'sh6a9b) : $signed(_GEN_10612); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10614 = 10'h175 == cnt[9:0] ? $signed(32'sh69e4) : $signed(_GEN_10613); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10615 = 10'h176 == cnt[9:0] ? $signed(32'sh692d) : $signed(_GEN_10614); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10616 = 10'h177 == cnt[9:0] ? $signed(32'sh6876) : $signed(_GEN_10615); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10617 = 10'h178 == cnt[9:0] ? $signed(32'sh67be) : $signed(_GEN_10616); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10618 = 10'h179 == cnt[9:0] ? $signed(32'sh6706) : $signed(_GEN_10617); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10619 = 10'h17a == cnt[9:0] ? $signed(32'sh664e) : $signed(_GEN_10618); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10620 = 10'h17b == cnt[9:0] ? $signed(32'sh6595) : $signed(_GEN_10619); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10621 = 10'h17c == cnt[9:0] ? $signed(32'sh64dd) : $signed(_GEN_10620); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10622 = 10'h17d == cnt[9:0] ? $signed(32'sh6424) : $signed(_GEN_10621); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10623 = 10'h17e == cnt[9:0] ? $signed(32'sh636b) : $signed(_GEN_10622); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10624 = 10'h17f == cnt[9:0] ? $signed(32'sh62b1) : $signed(_GEN_10623); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10625 = 10'h180 == cnt[9:0] ? $signed(32'sh61f8) : $signed(_GEN_10624); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10626 = 10'h181 == cnt[9:0] ? $signed(32'sh613e) : $signed(_GEN_10625); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10627 = 10'h182 == cnt[9:0] ? $signed(32'sh6084) : $signed(_GEN_10626); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10628 = 10'h183 == cnt[9:0] ? $signed(32'sh5fc9) : $signed(_GEN_10627); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10629 = 10'h184 == cnt[9:0] ? $signed(32'sh5f0f) : $signed(_GEN_10628); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10630 = 10'h185 == cnt[9:0] ? $signed(32'sh5e54) : $signed(_GEN_10629); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10631 = 10'h186 == cnt[9:0] ? $signed(32'sh5d99) : $signed(_GEN_10630); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10632 = 10'h187 == cnt[9:0] ? $signed(32'sh5cde) : $signed(_GEN_10631); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10633 = 10'h188 == cnt[9:0] ? $signed(32'sh5c22) : $signed(_GEN_10632); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10634 = 10'h189 == cnt[9:0] ? $signed(32'sh5b66) : $signed(_GEN_10633); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10635 = 10'h18a == cnt[9:0] ? $signed(32'sh5aaa) : $signed(_GEN_10634); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10636 = 10'h18b == cnt[9:0] ? $signed(32'sh59ee) : $signed(_GEN_10635); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10637 = 10'h18c == cnt[9:0] ? $signed(32'sh5932) : $signed(_GEN_10636); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10638 = 10'h18d == cnt[9:0] ? $signed(32'sh5875) : $signed(_GEN_10637); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10639 = 10'h18e == cnt[9:0] ? $signed(32'sh57b9) : $signed(_GEN_10638); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10640 = 10'h18f == cnt[9:0] ? $signed(32'sh56fc) : $signed(_GEN_10639); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10641 = 10'h190 == cnt[9:0] ? $signed(32'sh563e) : $signed(_GEN_10640); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10642 = 10'h191 == cnt[9:0] ? $signed(32'sh5581) : $signed(_GEN_10641); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10643 = 10'h192 == cnt[9:0] ? $signed(32'sh54c3) : $signed(_GEN_10642); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10644 = 10'h193 == cnt[9:0] ? $signed(32'sh5406) : $signed(_GEN_10643); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10645 = 10'h194 == cnt[9:0] ? $signed(32'sh5348) : $signed(_GEN_10644); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10646 = 10'h195 == cnt[9:0] ? $signed(32'sh5289) : $signed(_GEN_10645); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10647 = 10'h196 == cnt[9:0] ? $signed(32'sh51cb) : $signed(_GEN_10646); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10648 = 10'h197 == cnt[9:0] ? $signed(32'sh510c) : $signed(_GEN_10647); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10649 = 10'h198 == cnt[9:0] ? $signed(32'sh504d) : $signed(_GEN_10648); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10650 = 10'h199 == cnt[9:0] ? $signed(32'sh4f8e) : $signed(_GEN_10649); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10651 = 10'h19a == cnt[9:0] ? $signed(32'sh4ecf) : $signed(_GEN_10650); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10652 = 10'h19b == cnt[9:0] ? $signed(32'sh4e10) : $signed(_GEN_10651); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10653 = 10'h19c == cnt[9:0] ? $signed(32'sh4d50) : $signed(_GEN_10652); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10654 = 10'h19d == cnt[9:0] ? $signed(32'sh4c90) : $signed(_GEN_10653); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10655 = 10'h19e == cnt[9:0] ? $signed(32'sh4bd1) : $signed(_GEN_10654); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10656 = 10'h19f == cnt[9:0] ? $signed(32'sh4b10) : $signed(_GEN_10655); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10657 = 10'h1a0 == cnt[9:0] ? $signed(32'sh4a50) : $signed(_GEN_10656); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10658 = 10'h1a1 == cnt[9:0] ? $signed(32'sh4990) : $signed(_GEN_10657); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10659 = 10'h1a2 == cnt[9:0] ? $signed(32'sh48cf) : $signed(_GEN_10658); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10660 = 10'h1a3 == cnt[9:0] ? $signed(32'sh480e) : $signed(_GEN_10659); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10661 = 10'h1a4 == cnt[9:0] ? $signed(32'sh474d) : $signed(_GEN_10660); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10662 = 10'h1a5 == cnt[9:0] ? $signed(32'sh468c) : $signed(_GEN_10661); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10663 = 10'h1a6 == cnt[9:0] ? $signed(32'sh45cb) : $signed(_GEN_10662); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10664 = 10'h1a7 == cnt[9:0] ? $signed(32'sh4509) : $signed(_GEN_10663); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10665 = 10'h1a8 == cnt[9:0] ? $signed(32'sh4447) : $signed(_GEN_10664); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10666 = 10'h1a9 == cnt[9:0] ? $signed(32'sh4385) : $signed(_GEN_10665); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10667 = 10'h1aa == cnt[9:0] ? $signed(32'sh42c3) : $signed(_GEN_10666); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10668 = 10'h1ab == cnt[9:0] ? $signed(32'sh4201) : $signed(_GEN_10667); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10669 = 10'h1ac == cnt[9:0] ? $signed(32'sh413f) : $signed(_GEN_10668); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10670 = 10'h1ad == cnt[9:0] ? $signed(32'sh407c) : $signed(_GEN_10669); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10671 = 10'h1ae == cnt[9:0] ? $signed(32'sh3fba) : $signed(_GEN_10670); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10672 = 10'h1af == cnt[9:0] ? $signed(32'sh3ef7) : $signed(_GEN_10671); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10673 = 10'h1b0 == cnt[9:0] ? $signed(32'sh3e34) : $signed(_GEN_10672); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10674 = 10'h1b1 == cnt[9:0] ? $signed(32'sh3d71) : $signed(_GEN_10673); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10675 = 10'h1b2 == cnt[9:0] ? $signed(32'sh3cae) : $signed(_GEN_10674); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10676 = 10'h1b3 == cnt[9:0] ? $signed(32'sh3bea) : $signed(_GEN_10675); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10677 = 10'h1b4 == cnt[9:0] ? $signed(32'sh3b27) : $signed(_GEN_10676); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10678 = 10'h1b5 == cnt[9:0] ? $signed(32'sh3a63) : $signed(_GEN_10677); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10679 = 10'h1b6 == cnt[9:0] ? $signed(32'sh399f) : $signed(_GEN_10678); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10680 = 10'h1b7 == cnt[9:0] ? $signed(32'sh38db) : $signed(_GEN_10679); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10681 = 10'h1b8 == cnt[9:0] ? $signed(32'sh3817) : $signed(_GEN_10680); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10682 = 10'h1b9 == cnt[9:0] ? $signed(32'sh3753) : $signed(_GEN_10681); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10683 = 10'h1ba == cnt[9:0] ? $signed(32'sh368e) : $signed(_GEN_10682); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10684 = 10'h1bb == cnt[9:0] ? $signed(32'sh35ca) : $signed(_GEN_10683); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10685 = 10'h1bc == cnt[9:0] ? $signed(32'sh3505) : $signed(_GEN_10684); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10686 = 10'h1bd == cnt[9:0] ? $signed(32'sh3440) : $signed(_GEN_10685); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10687 = 10'h1be == cnt[9:0] ? $signed(32'sh337c) : $signed(_GEN_10686); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10688 = 10'h1bf == cnt[9:0] ? $signed(32'sh32b7) : $signed(_GEN_10687); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10689 = 10'h1c0 == cnt[9:0] ? $signed(32'sh31f1) : $signed(_GEN_10688); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10690 = 10'h1c1 == cnt[9:0] ? $signed(32'sh312c) : $signed(_GEN_10689); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10691 = 10'h1c2 == cnt[9:0] ? $signed(32'sh3067) : $signed(_GEN_10690); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10692 = 10'h1c3 == cnt[9:0] ? $signed(32'sh2fa1) : $signed(_GEN_10691); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10693 = 10'h1c4 == cnt[9:0] ? $signed(32'sh2edc) : $signed(_GEN_10692); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10694 = 10'h1c5 == cnt[9:0] ? $signed(32'sh2e16) : $signed(_GEN_10693); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10695 = 10'h1c6 == cnt[9:0] ? $signed(32'sh2d50) : $signed(_GEN_10694); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10696 = 10'h1c7 == cnt[9:0] ? $signed(32'sh2c8a) : $signed(_GEN_10695); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10697 = 10'h1c8 == cnt[9:0] ? $signed(32'sh2bc4) : $signed(_GEN_10696); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10698 = 10'h1c9 == cnt[9:0] ? $signed(32'sh2afe) : $signed(_GEN_10697); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10699 = 10'h1ca == cnt[9:0] ? $signed(32'sh2a38) : $signed(_GEN_10698); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10700 = 10'h1cb == cnt[9:0] ? $signed(32'sh2971) : $signed(_GEN_10699); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10701 = 10'h1cc == cnt[9:0] ? $signed(32'sh28ab) : $signed(_GEN_10700); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10702 = 10'h1cd == cnt[9:0] ? $signed(32'sh27e4) : $signed(_GEN_10701); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10703 = 10'h1ce == cnt[9:0] ? $signed(32'sh271e) : $signed(_GEN_10702); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10704 = 10'h1cf == cnt[9:0] ? $signed(32'sh2657) : $signed(_GEN_10703); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10705 = 10'h1d0 == cnt[9:0] ? $signed(32'sh2590) : $signed(_GEN_10704); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10706 = 10'h1d1 == cnt[9:0] ? $signed(32'sh24c9) : $signed(_GEN_10705); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10707 = 10'h1d2 == cnt[9:0] ? $signed(32'sh2402) : $signed(_GEN_10706); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10708 = 10'h1d3 == cnt[9:0] ? $signed(32'sh233b) : $signed(_GEN_10707); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10709 = 10'h1d4 == cnt[9:0] ? $signed(32'sh2274) : $signed(_GEN_10708); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10710 = 10'h1d5 == cnt[9:0] ? $signed(32'sh21ad) : $signed(_GEN_10709); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10711 = 10'h1d6 == cnt[9:0] ? $signed(32'sh20e5) : $signed(_GEN_10710); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10712 = 10'h1d7 == cnt[9:0] ? $signed(32'sh201e) : $signed(_GEN_10711); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10713 = 10'h1d8 == cnt[9:0] ? $signed(32'sh1f56) : $signed(_GEN_10712); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10714 = 10'h1d9 == cnt[9:0] ? $signed(32'sh1e8f) : $signed(_GEN_10713); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10715 = 10'h1da == cnt[9:0] ? $signed(32'sh1dc7) : $signed(_GEN_10714); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10716 = 10'h1db == cnt[9:0] ? $signed(32'sh1cff) : $signed(_GEN_10715); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10717 = 10'h1dc == cnt[9:0] ? $signed(32'sh1c38) : $signed(_GEN_10716); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10718 = 10'h1dd == cnt[9:0] ? $signed(32'sh1b70) : $signed(_GEN_10717); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10719 = 10'h1de == cnt[9:0] ? $signed(32'sh1aa8) : $signed(_GEN_10718); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10720 = 10'h1df == cnt[9:0] ? $signed(32'sh19e0) : $signed(_GEN_10719); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10721 = 10'h1e0 == cnt[9:0] ? $signed(32'sh1918) : $signed(_GEN_10720); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10722 = 10'h1e1 == cnt[9:0] ? $signed(32'sh1850) : $signed(_GEN_10721); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10723 = 10'h1e2 == cnt[9:0] ? $signed(32'sh1787) : $signed(_GEN_10722); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10724 = 10'h1e3 == cnt[9:0] ? $signed(32'sh16bf) : $signed(_GEN_10723); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10725 = 10'h1e4 == cnt[9:0] ? $signed(32'sh15f7) : $signed(_GEN_10724); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10726 = 10'h1e5 == cnt[9:0] ? $signed(32'sh152e) : $signed(_GEN_10725); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10727 = 10'h1e6 == cnt[9:0] ? $signed(32'sh1466) : $signed(_GEN_10726); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10728 = 10'h1e7 == cnt[9:0] ? $signed(32'sh139e) : $signed(_GEN_10727); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10729 = 10'h1e8 == cnt[9:0] ? $signed(32'sh12d5) : $signed(_GEN_10728); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10730 = 10'h1e9 == cnt[9:0] ? $signed(32'sh120d) : $signed(_GEN_10729); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10731 = 10'h1ea == cnt[9:0] ? $signed(32'sh1144) : $signed(_GEN_10730); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10732 = 10'h1eb == cnt[9:0] ? $signed(32'sh107b) : $signed(_GEN_10731); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10733 = 10'h1ec == cnt[9:0] ? $signed(32'shfb3) : $signed(_GEN_10732); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10734 = 10'h1ed == cnt[9:0] ? $signed(32'sheea) : $signed(_GEN_10733); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10735 = 10'h1ee == cnt[9:0] ? $signed(32'she21) : $signed(_GEN_10734); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10736 = 10'h1ef == cnt[9:0] ? $signed(32'shd59) : $signed(_GEN_10735); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10737 = 10'h1f0 == cnt[9:0] ? $signed(32'shc90) : $signed(_GEN_10736); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10738 = 10'h1f1 == cnt[9:0] ? $signed(32'shbc7) : $signed(_GEN_10737); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10739 = 10'h1f2 == cnt[9:0] ? $signed(32'shafe) : $signed(_GEN_10738); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10740 = 10'h1f3 == cnt[9:0] ? $signed(32'sha35) : $signed(_GEN_10739); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10741 = 10'h1f4 == cnt[9:0] ? $signed(32'sh96c) : $signed(_GEN_10740); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10742 = 10'h1f5 == cnt[9:0] ? $signed(32'sh8a3) : $signed(_GEN_10741); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10743 = 10'h1f6 == cnt[9:0] ? $signed(32'sh7da) : $signed(_GEN_10742); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10744 = 10'h1f7 == cnt[9:0] ? $signed(32'sh711) : $signed(_GEN_10743); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10745 = 10'h1f8 == cnt[9:0] ? $signed(32'sh648) : $signed(_GEN_10744); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10746 = 10'h1f9 == cnt[9:0] ? $signed(32'sh57f) : $signed(_GEN_10745); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10747 = 10'h1fa == cnt[9:0] ? $signed(32'sh4b6) : $signed(_GEN_10746); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10748 = 10'h1fb == cnt[9:0] ? $signed(32'sh3ed) : $signed(_GEN_10747); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10749 = 10'h1fc == cnt[9:0] ? $signed(32'sh324) : $signed(_GEN_10748); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10750 = 10'h1fd == cnt[9:0] ? $signed(32'sh25b) : $signed(_GEN_10749); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10751 = 10'h1fe == cnt[9:0] ? $signed(32'sh192) : $signed(_GEN_10750); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10752 = 10'h1ff == cnt[9:0] ? $signed(32'shc9) : $signed(_GEN_10751); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10753 = 10'h200 == cnt[9:0] ? $signed(32'sh0) : $signed(_GEN_10752); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10754 = 10'h201 == cnt[9:0] ? $signed(-32'shc9) : $signed(_GEN_10753); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10755 = 10'h202 == cnt[9:0] ? $signed(-32'sh192) : $signed(_GEN_10754); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10756 = 10'h203 == cnt[9:0] ? $signed(-32'sh25b) : $signed(_GEN_10755); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10757 = 10'h204 == cnt[9:0] ? $signed(-32'sh324) : $signed(_GEN_10756); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10758 = 10'h205 == cnt[9:0] ? $signed(-32'sh3ed) : $signed(_GEN_10757); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10759 = 10'h206 == cnt[9:0] ? $signed(-32'sh4b6) : $signed(_GEN_10758); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10760 = 10'h207 == cnt[9:0] ? $signed(-32'sh57f) : $signed(_GEN_10759); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10761 = 10'h208 == cnt[9:0] ? $signed(-32'sh648) : $signed(_GEN_10760); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10762 = 10'h209 == cnt[9:0] ? $signed(-32'sh711) : $signed(_GEN_10761); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10763 = 10'h20a == cnt[9:0] ? $signed(-32'sh7da) : $signed(_GEN_10762); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10764 = 10'h20b == cnt[9:0] ? $signed(-32'sh8a3) : $signed(_GEN_10763); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10765 = 10'h20c == cnt[9:0] ? $signed(-32'sh96c) : $signed(_GEN_10764); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10766 = 10'h20d == cnt[9:0] ? $signed(-32'sha35) : $signed(_GEN_10765); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10767 = 10'h20e == cnt[9:0] ? $signed(-32'shafe) : $signed(_GEN_10766); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10768 = 10'h20f == cnt[9:0] ? $signed(-32'shbc7) : $signed(_GEN_10767); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10769 = 10'h210 == cnt[9:0] ? $signed(-32'shc90) : $signed(_GEN_10768); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10770 = 10'h211 == cnt[9:0] ? $signed(-32'shd59) : $signed(_GEN_10769); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10771 = 10'h212 == cnt[9:0] ? $signed(-32'she21) : $signed(_GEN_10770); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10772 = 10'h213 == cnt[9:0] ? $signed(-32'sheea) : $signed(_GEN_10771); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10773 = 10'h214 == cnt[9:0] ? $signed(-32'shfb3) : $signed(_GEN_10772); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10774 = 10'h215 == cnt[9:0] ? $signed(-32'sh107b) : $signed(_GEN_10773); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10775 = 10'h216 == cnt[9:0] ? $signed(-32'sh1144) : $signed(_GEN_10774); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10776 = 10'h217 == cnt[9:0] ? $signed(-32'sh120d) : $signed(_GEN_10775); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10777 = 10'h218 == cnt[9:0] ? $signed(-32'sh12d5) : $signed(_GEN_10776); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10778 = 10'h219 == cnt[9:0] ? $signed(-32'sh139e) : $signed(_GEN_10777); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10779 = 10'h21a == cnt[9:0] ? $signed(-32'sh1466) : $signed(_GEN_10778); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10780 = 10'h21b == cnt[9:0] ? $signed(-32'sh152e) : $signed(_GEN_10779); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10781 = 10'h21c == cnt[9:0] ? $signed(-32'sh15f7) : $signed(_GEN_10780); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10782 = 10'h21d == cnt[9:0] ? $signed(-32'sh16bf) : $signed(_GEN_10781); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10783 = 10'h21e == cnt[9:0] ? $signed(-32'sh1787) : $signed(_GEN_10782); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10784 = 10'h21f == cnt[9:0] ? $signed(-32'sh1850) : $signed(_GEN_10783); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10785 = 10'h220 == cnt[9:0] ? $signed(-32'sh1918) : $signed(_GEN_10784); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10786 = 10'h221 == cnt[9:0] ? $signed(-32'sh19e0) : $signed(_GEN_10785); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10787 = 10'h222 == cnt[9:0] ? $signed(-32'sh1aa8) : $signed(_GEN_10786); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10788 = 10'h223 == cnt[9:0] ? $signed(-32'sh1b70) : $signed(_GEN_10787); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10789 = 10'h224 == cnt[9:0] ? $signed(-32'sh1c38) : $signed(_GEN_10788); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10790 = 10'h225 == cnt[9:0] ? $signed(-32'sh1cff) : $signed(_GEN_10789); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10791 = 10'h226 == cnt[9:0] ? $signed(-32'sh1dc7) : $signed(_GEN_10790); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10792 = 10'h227 == cnt[9:0] ? $signed(-32'sh1e8f) : $signed(_GEN_10791); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10793 = 10'h228 == cnt[9:0] ? $signed(-32'sh1f56) : $signed(_GEN_10792); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10794 = 10'h229 == cnt[9:0] ? $signed(-32'sh201e) : $signed(_GEN_10793); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10795 = 10'h22a == cnt[9:0] ? $signed(-32'sh20e5) : $signed(_GEN_10794); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10796 = 10'h22b == cnt[9:0] ? $signed(-32'sh21ad) : $signed(_GEN_10795); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10797 = 10'h22c == cnt[9:0] ? $signed(-32'sh2274) : $signed(_GEN_10796); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10798 = 10'h22d == cnt[9:0] ? $signed(-32'sh233b) : $signed(_GEN_10797); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10799 = 10'h22e == cnt[9:0] ? $signed(-32'sh2402) : $signed(_GEN_10798); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10800 = 10'h22f == cnt[9:0] ? $signed(-32'sh24c9) : $signed(_GEN_10799); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10801 = 10'h230 == cnt[9:0] ? $signed(-32'sh2590) : $signed(_GEN_10800); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10802 = 10'h231 == cnt[9:0] ? $signed(-32'sh2657) : $signed(_GEN_10801); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10803 = 10'h232 == cnt[9:0] ? $signed(-32'sh271e) : $signed(_GEN_10802); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10804 = 10'h233 == cnt[9:0] ? $signed(-32'sh27e4) : $signed(_GEN_10803); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10805 = 10'h234 == cnt[9:0] ? $signed(-32'sh28ab) : $signed(_GEN_10804); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10806 = 10'h235 == cnt[9:0] ? $signed(-32'sh2971) : $signed(_GEN_10805); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10807 = 10'h236 == cnt[9:0] ? $signed(-32'sh2a38) : $signed(_GEN_10806); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10808 = 10'h237 == cnt[9:0] ? $signed(-32'sh2afe) : $signed(_GEN_10807); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10809 = 10'h238 == cnt[9:0] ? $signed(-32'sh2bc4) : $signed(_GEN_10808); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10810 = 10'h239 == cnt[9:0] ? $signed(-32'sh2c8a) : $signed(_GEN_10809); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10811 = 10'h23a == cnt[9:0] ? $signed(-32'sh2d50) : $signed(_GEN_10810); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10812 = 10'h23b == cnt[9:0] ? $signed(-32'sh2e16) : $signed(_GEN_10811); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10813 = 10'h23c == cnt[9:0] ? $signed(-32'sh2edc) : $signed(_GEN_10812); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10814 = 10'h23d == cnt[9:0] ? $signed(-32'sh2fa1) : $signed(_GEN_10813); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10815 = 10'h23e == cnt[9:0] ? $signed(-32'sh3067) : $signed(_GEN_10814); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10816 = 10'h23f == cnt[9:0] ? $signed(-32'sh312c) : $signed(_GEN_10815); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10817 = 10'h240 == cnt[9:0] ? $signed(-32'sh31f1) : $signed(_GEN_10816); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10818 = 10'h241 == cnt[9:0] ? $signed(-32'sh32b7) : $signed(_GEN_10817); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10819 = 10'h242 == cnt[9:0] ? $signed(-32'sh337c) : $signed(_GEN_10818); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10820 = 10'h243 == cnt[9:0] ? $signed(-32'sh3440) : $signed(_GEN_10819); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10821 = 10'h244 == cnt[9:0] ? $signed(-32'sh3505) : $signed(_GEN_10820); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10822 = 10'h245 == cnt[9:0] ? $signed(-32'sh35ca) : $signed(_GEN_10821); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10823 = 10'h246 == cnt[9:0] ? $signed(-32'sh368e) : $signed(_GEN_10822); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10824 = 10'h247 == cnt[9:0] ? $signed(-32'sh3753) : $signed(_GEN_10823); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10825 = 10'h248 == cnt[9:0] ? $signed(-32'sh3817) : $signed(_GEN_10824); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10826 = 10'h249 == cnt[9:0] ? $signed(-32'sh38db) : $signed(_GEN_10825); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10827 = 10'h24a == cnt[9:0] ? $signed(-32'sh399f) : $signed(_GEN_10826); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10828 = 10'h24b == cnt[9:0] ? $signed(-32'sh3a63) : $signed(_GEN_10827); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10829 = 10'h24c == cnt[9:0] ? $signed(-32'sh3b27) : $signed(_GEN_10828); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10830 = 10'h24d == cnt[9:0] ? $signed(-32'sh3bea) : $signed(_GEN_10829); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10831 = 10'h24e == cnt[9:0] ? $signed(-32'sh3cae) : $signed(_GEN_10830); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10832 = 10'h24f == cnt[9:0] ? $signed(-32'sh3d71) : $signed(_GEN_10831); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10833 = 10'h250 == cnt[9:0] ? $signed(-32'sh3e34) : $signed(_GEN_10832); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10834 = 10'h251 == cnt[9:0] ? $signed(-32'sh3ef7) : $signed(_GEN_10833); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10835 = 10'h252 == cnt[9:0] ? $signed(-32'sh3fba) : $signed(_GEN_10834); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10836 = 10'h253 == cnt[9:0] ? $signed(-32'sh407c) : $signed(_GEN_10835); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10837 = 10'h254 == cnt[9:0] ? $signed(-32'sh413f) : $signed(_GEN_10836); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10838 = 10'h255 == cnt[9:0] ? $signed(-32'sh4201) : $signed(_GEN_10837); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10839 = 10'h256 == cnt[9:0] ? $signed(-32'sh42c3) : $signed(_GEN_10838); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10840 = 10'h257 == cnt[9:0] ? $signed(-32'sh4385) : $signed(_GEN_10839); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10841 = 10'h258 == cnt[9:0] ? $signed(-32'sh4447) : $signed(_GEN_10840); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10842 = 10'h259 == cnt[9:0] ? $signed(-32'sh4509) : $signed(_GEN_10841); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10843 = 10'h25a == cnt[9:0] ? $signed(-32'sh45cb) : $signed(_GEN_10842); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10844 = 10'h25b == cnt[9:0] ? $signed(-32'sh468c) : $signed(_GEN_10843); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10845 = 10'h25c == cnt[9:0] ? $signed(-32'sh474d) : $signed(_GEN_10844); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10846 = 10'h25d == cnt[9:0] ? $signed(-32'sh480e) : $signed(_GEN_10845); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10847 = 10'h25e == cnt[9:0] ? $signed(-32'sh48cf) : $signed(_GEN_10846); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10848 = 10'h25f == cnt[9:0] ? $signed(-32'sh4990) : $signed(_GEN_10847); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10849 = 10'h260 == cnt[9:0] ? $signed(-32'sh4a50) : $signed(_GEN_10848); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10850 = 10'h261 == cnt[9:0] ? $signed(-32'sh4b10) : $signed(_GEN_10849); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10851 = 10'h262 == cnt[9:0] ? $signed(-32'sh4bd1) : $signed(_GEN_10850); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10852 = 10'h263 == cnt[9:0] ? $signed(-32'sh4c90) : $signed(_GEN_10851); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10853 = 10'h264 == cnt[9:0] ? $signed(-32'sh4d50) : $signed(_GEN_10852); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10854 = 10'h265 == cnt[9:0] ? $signed(-32'sh4e10) : $signed(_GEN_10853); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10855 = 10'h266 == cnt[9:0] ? $signed(-32'sh4ecf) : $signed(_GEN_10854); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10856 = 10'h267 == cnt[9:0] ? $signed(-32'sh4f8e) : $signed(_GEN_10855); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10857 = 10'h268 == cnt[9:0] ? $signed(-32'sh504d) : $signed(_GEN_10856); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10858 = 10'h269 == cnt[9:0] ? $signed(-32'sh510c) : $signed(_GEN_10857); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10859 = 10'h26a == cnt[9:0] ? $signed(-32'sh51cb) : $signed(_GEN_10858); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10860 = 10'h26b == cnt[9:0] ? $signed(-32'sh5289) : $signed(_GEN_10859); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10861 = 10'h26c == cnt[9:0] ? $signed(-32'sh5348) : $signed(_GEN_10860); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10862 = 10'h26d == cnt[9:0] ? $signed(-32'sh5406) : $signed(_GEN_10861); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10863 = 10'h26e == cnt[9:0] ? $signed(-32'sh54c3) : $signed(_GEN_10862); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10864 = 10'h26f == cnt[9:0] ? $signed(-32'sh5581) : $signed(_GEN_10863); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10865 = 10'h270 == cnt[9:0] ? $signed(-32'sh563e) : $signed(_GEN_10864); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10866 = 10'h271 == cnt[9:0] ? $signed(-32'sh56fc) : $signed(_GEN_10865); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10867 = 10'h272 == cnt[9:0] ? $signed(-32'sh57b9) : $signed(_GEN_10866); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10868 = 10'h273 == cnt[9:0] ? $signed(-32'sh5875) : $signed(_GEN_10867); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10869 = 10'h274 == cnt[9:0] ? $signed(-32'sh5932) : $signed(_GEN_10868); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10870 = 10'h275 == cnt[9:0] ? $signed(-32'sh59ee) : $signed(_GEN_10869); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10871 = 10'h276 == cnt[9:0] ? $signed(-32'sh5aaa) : $signed(_GEN_10870); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10872 = 10'h277 == cnt[9:0] ? $signed(-32'sh5b66) : $signed(_GEN_10871); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10873 = 10'h278 == cnt[9:0] ? $signed(-32'sh5c22) : $signed(_GEN_10872); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10874 = 10'h279 == cnt[9:0] ? $signed(-32'sh5cde) : $signed(_GEN_10873); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10875 = 10'h27a == cnt[9:0] ? $signed(-32'sh5d99) : $signed(_GEN_10874); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10876 = 10'h27b == cnt[9:0] ? $signed(-32'sh5e54) : $signed(_GEN_10875); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10877 = 10'h27c == cnt[9:0] ? $signed(-32'sh5f0f) : $signed(_GEN_10876); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10878 = 10'h27d == cnt[9:0] ? $signed(-32'sh5fc9) : $signed(_GEN_10877); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10879 = 10'h27e == cnt[9:0] ? $signed(-32'sh6084) : $signed(_GEN_10878); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10880 = 10'h27f == cnt[9:0] ? $signed(-32'sh613e) : $signed(_GEN_10879); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10881 = 10'h280 == cnt[9:0] ? $signed(-32'sh61f8) : $signed(_GEN_10880); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10882 = 10'h281 == cnt[9:0] ? $signed(-32'sh62b1) : $signed(_GEN_10881); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10883 = 10'h282 == cnt[9:0] ? $signed(-32'sh636b) : $signed(_GEN_10882); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10884 = 10'h283 == cnt[9:0] ? $signed(-32'sh6424) : $signed(_GEN_10883); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10885 = 10'h284 == cnt[9:0] ? $signed(-32'sh64dd) : $signed(_GEN_10884); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10886 = 10'h285 == cnt[9:0] ? $signed(-32'sh6595) : $signed(_GEN_10885); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10887 = 10'h286 == cnt[9:0] ? $signed(-32'sh664e) : $signed(_GEN_10886); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10888 = 10'h287 == cnt[9:0] ? $signed(-32'sh6706) : $signed(_GEN_10887); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10889 = 10'h288 == cnt[9:0] ? $signed(-32'sh67be) : $signed(_GEN_10888); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10890 = 10'h289 == cnt[9:0] ? $signed(-32'sh6876) : $signed(_GEN_10889); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10891 = 10'h28a == cnt[9:0] ? $signed(-32'sh692d) : $signed(_GEN_10890); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10892 = 10'h28b == cnt[9:0] ? $signed(-32'sh69e4) : $signed(_GEN_10891); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10893 = 10'h28c == cnt[9:0] ? $signed(-32'sh6a9b) : $signed(_GEN_10892); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10894 = 10'h28d == cnt[9:0] ? $signed(-32'sh6b52) : $signed(_GEN_10893); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10895 = 10'h28e == cnt[9:0] ? $signed(-32'sh6c08) : $signed(_GEN_10894); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10896 = 10'h28f == cnt[9:0] ? $signed(-32'sh6cbe) : $signed(_GEN_10895); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10897 = 10'h290 == cnt[9:0] ? $signed(-32'sh6d74) : $signed(_GEN_10896); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10898 = 10'h291 == cnt[9:0] ? $signed(-32'sh6e2a) : $signed(_GEN_10897); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10899 = 10'h292 == cnt[9:0] ? $signed(-32'sh6edf) : $signed(_GEN_10898); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10900 = 10'h293 == cnt[9:0] ? $signed(-32'sh6f94) : $signed(_GEN_10899); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10901 = 10'h294 == cnt[9:0] ? $signed(-32'sh7049) : $signed(_GEN_10900); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10902 = 10'h295 == cnt[9:0] ? $signed(-32'sh70fe) : $signed(_GEN_10901); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10903 = 10'h296 == cnt[9:0] ? $signed(-32'sh71b2) : $signed(_GEN_10902); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10904 = 10'h297 == cnt[9:0] ? $signed(-32'sh7266) : $signed(_GEN_10903); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10905 = 10'h298 == cnt[9:0] ? $signed(-32'sh731a) : $signed(_GEN_10904); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10906 = 10'h299 == cnt[9:0] ? $signed(-32'sh73cd) : $signed(_GEN_10905); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10907 = 10'h29a == cnt[9:0] ? $signed(-32'sh7480) : $signed(_GEN_10906); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10908 = 10'h29b == cnt[9:0] ? $signed(-32'sh7533) : $signed(_GEN_10907); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10909 = 10'h29c == cnt[9:0] ? $signed(-32'sh75e6) : $signed(_GEN_10908); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10910 = 10'h29d == cnt[9:0] ? $signed(-32'sh7698) : $signed(_GEN_10909); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10911 = 10'h29e == cnt[9:0] ? $signed(-32'sh774a) : $signed(_GEN_10910); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10912 = 10'h29f == cnt[9:0] ? $signed(-32'sh77fc) : $signed(_GEN_10911); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10913 = 10'h2a0 == cnt[9:0] ? $signed(-32'sh78ad) : $signed(_GEN_10912); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10914 = 10'h2a1 == cnt[9:0] ? $signed(-32'sh795f) : $signed(_GEN_10913); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10915 = 10'h2a2 == cnt[9:0] ? $signed(-32'sh7a10) : $signed(_GEN_10914); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10916 = 10'h2a3 == cnt[9:0] ? $signed(-32'sh7ac0) : $signed(_GEN_10915); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10917 = 10'h2a4 == cnt[9:0] ? $signed(-32'sh7b70) : $signed(_GEN_10916); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10918 = 10'h2a5 == cnt[9:0] ? $signed(-32'sh7c20) : $signed(_GEN_10917); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10919 = 10'h2a6 == cnt[9:0] ? $signed(-32'sh7cd0) : $signed(_GEN_10918); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10920 = 10'h2a7 == cnt[9:0] ? $signed(-32'sh7d7f) : $signed(_GEN_10919); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10921 = 10'h2a8 == cnt[9:0] ? $signed(-32'sh7e2f) : $signed(_GEN_10920); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10922 = 10'h2a9 == cnt[9:0] ? $signed(-32'sh7edd) : $signed(_GEN_10921); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10923 = 10'h2aa == cnt[9:0] ? $signed(-32'sh7f8c) : $signed(_GEN_10922); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10924 = 10'h2ab == cnt[9:0] ? $signed(-32'sh803a) : $signed(_GEN_10923); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10925 = 10'h2ac == cnt[9:0] ? $signed(-32'sh80e8) : $signed(_GEN_10924); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10926 = 10'h2ad == cnt[9:0] ? $signed(-32'sh8195) : $signed(_GEN_10925); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10927 = 10'h2ae == cnt[9:0] ? $signed(-32'sh8243) : $signed(_GEN_10926); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10928 = 10'h2af == cnt[9:0] ? $signed(-32'sh82f0) : $signed(_GEN_10927); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10929 = 10'h2b0 == cnt[9:0] ? $signed(-32'sh839c) : $signed(_GEN_10928); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10930 = 10'h2b1 == cnt[9:0] ? $signed(-32'sh8449) : $signed(_GEN_10929); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10931 = 10'h2b2 == cnt[9:0] ? $signed(-32'sh84f5) : $signed(_GEN_10930); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10932 = 10'h2b3 == cnt[9:0] ? $signed(-32'sh85a0) : $signed(_GEN_10931); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10933 = 10'h2b4 == cnt[9:0] ? $signed(-32'sh864c) : $signed(_GEN_10932); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10934 = 10'h2b5 == cnt[9:0] ? $signed(-32'sh86f7) : $signed(_GEN_10933); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10935 = 10'h2b6 == cnt[9:0] ? $signed(-32'sh87a1) : $signed(_GEN_10934); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10936 = 10'h2b7 == cnt[9:0] ? $signed(-32'sh884c) : $signed(_GEN_10935); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10937 = 10'h2b8 == cnt[9:0] ? $signed(-32'sh88f6) : $signed(_GEN_10936); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10938 = 10'h2b9 == cnt[9:0] ? $signed(-32'sh899f) : $signed(_GEN_10937); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10939 = 10'h2ba == cnt[9:0] ? $signed(-32'sh8a49) : $signed(_GEN_10938); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10940 = 10'h2bb == cnt[9:0] ? $signed(-32'sh8af2) : $signed(_GEN_10939); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10941 = 10'h2bc == cnt[9:0] ? $signed(-32'sh8b9a) : $signed(_GEN_10940); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10942 = 10'h2bd == cnt[9:0] ? $signed(-32'sh8c43) : $signed(_GEN_10941); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10943 = 10'h2be == cnt[9:0] ? $signed(-32'sh8ceb) : $signed(_GEN_10942); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10944 = 10'h2bf == cnt[9:0] ? $signed(-32'sh8d93) : $signed(_GEN_10943); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10945 = 10'h2c0 == cnt[9:0] ? $signed(-32'sh8e3a) : $signed(_GEN_10944); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10946 = 10'h2c1 == cnt[9:0] ? $signed(-32'sh8ee1) : $signed(_GEN_10945); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10947 = 10'h2c2 == cnt[9:0] ? $signed(-32'sh8f88) : $signed(_GEN_10946); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10948 = 10'h2c3 == cnt[9:0] ? $signed(-32'sh902e) : $signed(_GEN_10947); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10949 = 10'h2c4 == cnt[9:0] ? $signed(-32'sh90d4) : $signed(_GEN_10948); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10950 = 10'h2c5 == cnt[9:0] ? $signed(-32'sh9179) : $signed(_GEN_10949); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10951 = 10'h2c6 == cnt[9:0] ? $signed(-32'sh921f) : $signed(_GEN_10950); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10952 = 10'h2c7 == cnt[9:0] ? $signed(-32'sh92c4) : $signed(_GEN_10951); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10953 = 10'h2c8 == cnt[9:0] ? $signed(-32'sh9368) : $signed(_GEN_10952); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10954 = 10'h2c9 == cnt[9:0] ? $signed(-32'sh940c) : $signed(_GEN_10953); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10955 = 10'h2ca == cnt[9:0] ? $signed(-32'sh94b0) : $signed(_GEN_10954); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10956 = 10'h2cb == cnt[9:0] ? $signed(-32'sh9554) : $signed(_GEN_10955); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10957 = 10'h2cc == cnt[9:0] ? $signed(-32'sh95f7) : $signed(_GEN_10956); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10958 = 10'h2cd == cnt[9:0] ? $signed(-32'sh969a) : $signed(_GEN_10957); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10959 = 10'h2ce == cnt[9:0] ? $signed(-32'sh973c) : $signed(_GEN_10958); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10960 = 10'h2cf == cnt[9:0] ? $signed(-32'sh97de) : $signed(_GEN_10959); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10961 = 10'h2d0 == cnt[9:0] ? $signed(-32'sh9880) : $signed(_GEN_10960); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10962 = 10'h2d1 == cnt[9:0] ? $signed(-32'sh9921) : $signed(_GEN_10961); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10963 = 10'h2d2 == cnt[9:0] ? $signed(-32'sh99c2) : $signed(_GEN_10962); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10964 = 10'h2d3 == cnt[9:0] ? $signed(-32'sh9a63) : $signed(_GEN_10963); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10965 = 10'h2d4 == cnt[9:0] ? $signed(-32'sh9b03) : $signed(_GEN_10964); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10966 = 10'h2d5 == cnt[9:0] ? $signed(-32'sh9ba3) : $signed(_GEN_10965); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10967 = 10'h2d6 == cnt[9:0] ? $signed(-32'sh9c42) : $signed(_GEN_10966); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10968 = 10'h2d7 == cnt[9:0] ? $signed(-32'sh9ce1) : $signed(_GEN_10967); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10969 = 10'h2d8 == cnt[9:0] ? $signed(-32'sh9d80) : $signed(_GEN_10968); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10970 = 10'h2d9 == cnt[9:0] ? $signed(-32'sh9e1e) : $signed(_GEN_10969); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10971 = 10'h2da == cnt[9:0] ? $signed(-32'sh9ebc) : $signed(_GEN_10970); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10972 = 10'h2db == cnt[9:0] ? $signed(-32'sh9f5a) : $signed(_GEN_10971); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10973 = 10'h2dc == cnt[9:0] ? $signed(-32'sh9ff7) : $signed(_GEN_10972); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10974 = 10'h2dd == cnt[9:0] ? $signed(-32'sha094) : $signed(_GEN_10973); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10975 = 10'h2de == cnt[9:0] ? $signed(-32'sha130) : $signed(_GEN_10974); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10976 = 10'h2df == cnt[9:0] ? $signed(-32'sha1cc) : $signed(_GEN_10975); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10977 = 10'h2e0 == cnt[9:0] ? $signed(-32'sha268) : $signed(_GEN_10976); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10978 = 10'h2e1 == cnt[9:0] ? $signed(-32'sha303) : $signed(_GEN_10977); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10979 = 10'h2e2 == cnt[9:0] ? $signed(-32'sha39e) : $signed(_GEN_10978); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10980 = 10'h2e3 == cnt[9:0] ? $signed(-32'sha438) : $signed(_GEN_10979); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10981 = 10'h2e4 == cnt[9:0] ? $signed(-32'sha4d2) : $signed(_GEN_10980); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10982 = 10'h2e5 == cnt[9:0] ? $signed(-32'sha56c) : $signed(_GEN_10981); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10983 = 10'h2e6 == cnt[9:0] ? $signed(-32'sha605) : $signed(_GEN_10982); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10984 = 10'h2e7 == cnt[9:0] ? $signed(-32'sha69e) : $signed(_GEN_10983); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10985 = 10'h2e8 == cnt[9:0] ? $signed(-32'sha736) : $signed(_GEN_10984); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10986 = 10'h2e9 == cnt[9:0] ? $signed(-32'sha7ce) : $signed(_GEN_10985); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10987 = 10'h2ea == cnt[9:0] ? $signed(-32'sha866) : $signed(_GEN_10986); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10988 = 10'h2eb == cnt[9:0] ? $signed(-32'sha8fd) : $signed(_GEN_10987); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10989 = 10'h2ec == cnt[9:0] ? $signed(-32'sha994) : $signed(_GEN_10988); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10990 = 10'h2ed == cnt[9:0] ? $signed(-32'shaa2a) : $signed(_GEN_10989); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10991 = 10'h2ee == cnt[9:0] ? $signed(-32'shaac1) : $signed(_GEN_10990); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10992 = 10'h2ef == cnt[9:0] ? $signed(-32'shab56) : $signed(_GEN_10991); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10993 = 10'h2f0 == cnt[9:0] ? $signed(-32'shabeb) : $signed(_GEN_10992); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10994 = 10'h2f1 == cnt[9:0] ? $signed(-32'shac80) : $signed(_GEN_10993); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10995 = 10'h2f2 == cnt[9:0] ? $signed(-32'shad14) : $signed(_GEN_10994); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10996 = 10'h2f3 == cnt[9:0] ? $signed(-32'shada8) : $signed(_GEN_10995); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10997 = 10'h2f4 == cnt[9:0] ? $signed(-32'shae3c) : $signed(_GEN_10996); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10998 = 10'h2f5 == cnt[9:0] ? $signed(-32'shaecf) : $signed(_GEN_10997); // @[FFT.scala 34:12]
  wire [31:0] _GEN_10999 = 10'h2f6 == cnt[9:0] ? $signed(-32'shaf62) : $signed(_GEN_10998); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11000 = 10'h2f7 == cnt[9:0] ? $signed(-32'shaff4) : $signed(_GEN_10999); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11001 = 10'h2f8 == cnt[9:0] ? $signed(-32'shb086) : $signed(_GEN_11000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11002 = 10'h2f9 == cnt[9:0] ? $signed(-32'shb117) : $signed(_GEN_11001); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11003 = 10'h2fa == cnt[9:0] ? $signed(-32'shb1a8) : $signed(_GEN_11002); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11004 = 10'h2fb == cnt[9:0] ? $signed(-32'shb239) : $signed(_GEN_11003); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11005 = 10'h2fc == cnt[9:0] ? $signed(-32'shb2c9) : $signed(_GEN_11004); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11006 = 10'h2fd == cnt[9:0] ? $signed(-32'shb358) : $signed(_GEN_11005); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11007 = 10'h2fe == cnt[9:0] ? $signed(-32'shb3e8) : $signed(_GEN_11006); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11008 = 10'h2ff == cnt[9:0] ? $signed(-32'shb477) : $signed(_GEN_11007); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11009 = 10'h300 == cnt[9:0] ? $signed(-32'shb505) : $signed(_GEN_11008); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11010 = 10'h301 == cnt[9:0] ? $signed(-32'shb593) : $signed(_GEN_11009); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11011 = 10'h302 == cnt[9:0] ? $signed(-32'shb620) : $signed(_GEN_11010); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11012 = 10'h303 == cnt[9:0] ? $signed(-32'shb6ad) : $signed(_GEN_11011); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11013 = 10'h304 == cnt[9:0] ? $signed(-32'shb73a) : $signed(_GEN_11012); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11014 = 10'h305 == cnt[9:0] ? $signed(-32'shb7c6) : $signed(_GEN_11013); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11015 = 10'h306 == cnt[9:0] ? $signed(-32'shb852) : $signed(_GEN_11014); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11016 = 10'h307 == cnt[9:0] ? $signed(-32'shb8dd) : $signed(_GEN_11015); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11017 = 10'h308 == cnt[9:0] ? $signed(-32'shb968) : $signed(_GEN_11016); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11018 = 10'h309 == cnt[9:0] ? $signed(-32'shb9f3) : $signed(_GEN_11017); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11019 = 10'h30a == cnt[9:0] ? $signed(-32'shba7d) : $signed(_GEN_11018); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11020 = 10'h30b == cnt[9:0] ? $signed(-32'shbb06) : $signed(_GEN_11019); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11021 = 10'h30c == cnt[9:0] ? $signed(-32'shbb8f) : $signed(_GEN_11020); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11022 = 10'h30d == cnt[9:0] ? $signed(-32'shbc18) : $signed(_GEN_11021); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11023 = 10'h30e == cnt[9:0] ? $signed(-32'shbca0) : $signed(_GEN_11022); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11024 = 10'h30f == cnt[9:0] ? $signed(-32'shbd28) : $signed(_GEN_11023); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11025 = 10'h310 == cnt[9:0] ? $signed(-32'shbdaf) : $signed(_GEN_11024); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11026 = 10'h311 == cnt[9:0] ? $signed(-32'shbe36) : $signed(_GEN_11025); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11027 = 10'h312 == cnt[9:0] ? $signed(-32'shbebc) : $signed(_GEN_11026); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11028 = 10'h313 == cnt[9:0] ? $signed(-32'shbf42) : $signed(_GEN_11027); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11029 = 10'h314 == cnt[9:0] ? $signed(-32'shbfc7) : $signed(_GEN_11028); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11030 = 10'h315 == cnt[9:0] ? $signed(-32'shc04c) : $signed(_GEN_11029); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11031 = 10'h316 == cnt[9:0] ? $signed(-32'shc0d1) : $signed(_GEN_11030); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11032 = 10'h317 == cnt[9:0] ? $signed(-32'shc155) : $signed(_GEN_11031); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11033 = 10'h318 == cnt[9:0] ? $signed(-32'shc1d8) : $signed(_GEN_11032); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11034 = 10'h319 == cnt[9:0] ? $signed(-32'shc25c) : $signed(_GEN_11033); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11035 = 10'h31a == cnt[9:0] ? $signed(-32'shc2de) : $signed(_GEN_11034); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11036 = 10'h31b == cnt[9:0] ? $signed(-32'shc360) : $signed(_GEN_11035); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11037 = 10'h31c == cnt[9:0] ? $signed(-32'shc3e2) : $signed(_GEN_11036); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11038 = 10'h31d == cnt[9:0] ? $signed(-32'shc463) : $signed(_GEN_11037); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11039 = 10'h31e == cnt[9:0] ? $signed(-32'shc4e4) : $signed(_GEN_11038); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11040 = 10'h31f == cnt[9:0] ? $signed(-32'shc564) : $signed(_GEN_11039); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11041 = 10'h320 == cnt[9:0] ? $signed(-32'shc5e4) : $signed(_GEN_11040); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11042 = 10'h321 == cnt[9:0] ? $signed(-32'shc663) : $signed(_GEN_11041); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11043 = 10'h322 == cnt[9:0] ? $signed(-32'shc6e2) : $signed(_GEN_11042); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11044 = 10'h323 == cnt[9:0] ? $signed(-32'shc761) : $signed(_GEN_11043); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11045 = 10'h324 == cnt[9:0] ? $signed(-32'shc7de) : $signed(_GEN_11044); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11046 = 10'h325 == cnt[9:0] ? $signed(-32'shc85c) : $signed(_GEN_11045); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11047 = 10'h326 == cnt[9:0] ? $signed(-32'shc8d9) : $signed(_GEN_11046); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11048 = 10'h327 == cnt[9:0] ? $signed(-32'shc955) : $signed(_GEN_11047); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11049 = 10'h328 == cnt[9:0] ? $signed(-32'shc9d1) : $signed(_GEN_11048); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11050 = 10'h329 == cnt[9:0] ? $signed(-32'shca4d) : $signed(_GEN_11049); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11051 = 10'h32a == cnt[9:0] ? $signed(-32'shcac7) : $signed(_GEN_11050); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11052 = 10'h32b == cnt[9:0] ? $signed(-32'shcb42) : $signed(_GEN_11051); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11053 = 10'h32c == cnt[9:0] ? $signed(-32'shcbbc) : $signed(_GEN_11052); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11054 = 10'h32d == cnt[9:0] ? $signed(-32'shcc35) : $signed(_GEN_11053); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11055 = 10'h32e == cnt[9:0] ? $signed(-32'shccae) : $signed(_GEN_11054); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11056 = 10'h32f == cnt[9:0] ? $signed(-32'shcd27) : $signed(_GEN_11055); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11057 = 10'h330 == cnt[9:0] ? $signed(-32'shcd9f) : $signed(_GEN_11056); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11058 = 10'h331 == cnt[9:0] ? $signed(-32'shce17) : $signed(_GEN_11057); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11059 = 10'h332 == cnt[9:0] ? $signed(-32'shce8e) : $signed(_GEN_11058); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11060 = 10'h333 == cnt[9:0] ? $signed(-32'shcf04) : $signed(_GEN_11059); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11061 = 10'h334 == cnt[9:0] ? $signed(-32'shcf7a) : $signed(_GEN_11060); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11062 = 10'h335 == cnt[9:0] ? $signed(-32'shcff0) : $signed(_GEN_11061); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11063 = 10'h336 == cnt[9:0] ? $signed(-32'shd065) : $signed(_GEN_11062); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11064 = 10'h337 == cnt[9:0] ? $signed(-32'shd0d9) : $signed(_GEN_11063); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11065 = 10'h338 == cnt[9:0] ? $signed(-32'shd14d) : $signed(_GEN_11064); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11066 = 10'h339 == cnt[9:0] ? $signed(-32'shd1c1) : $signed(_GEN_11065); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11067 = 10'h33a == cnt[9:0] ? $signed(-32'shd234) : $signed(_GEN_11066); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11068 = 10'h33b == cnt[9:0] ? $signed(-32'shd2a6) : $signed(_GEN_11067); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11069 = 10'h33c == cnt[9:0] ? $signed(-32'shd318) : $signed(_GEN_11068); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11070 = 10'h33d == cnt[9:0] ? $signed(-32'shd38a) : $signed(_GEN_11069); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11071 = 10'h33e == cnt[9:0] ? $signed(-32'shd3fb) : $signed(_GEN_11070); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11072 = 10'h33f == cnt[9:0] ? $signed(-32'shd46b) : $signed(_GEN_11071); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11073 = 10'h340 == cnt[9:0] ? $signed(-32'shd4db) : $signed(_GEN_11072); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11074 = 10'h341 == cnt[9:0] ? $signed(-32'shd54b) : $signed(_GEN_11073); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11075 = 10'h342 == cnt[9:0] ? $signed(-32'shd5ba) : $signed(_GEN_11074); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11076 = 10'h343 == cnt[9:0] ? $signed(-32'shd628) : $signed(_GEN_11075); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11077 = 10'h344 == cnt[9:0] ? $signed(-32'shd696) : $signed(_GEN_11076); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11078 = 10'h345 == cnt[9:0] ? $signed(-32'shd703) : $signed(_GEN_11077); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11079 = 10'h346 == cnt[9:0] ? $signed(-32'shd770) : $signed(_GEN_11078); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11080 = 10'h347 == cnt[9:0] ? $signed(-32'shd7dc) : $signed(_GEN_11079); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11081 = 10'h348 == cnt[9:0] ? $signed(-32'shd848) : $signed(_GEN_11080); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11082 = 10'h349 == cnt[9:0] ? $signed(-32'shd8b4) : $signed(_GEN_11081); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11083 = 10'h34a == cnt[9:0] ? $signed(-32'shd91e) : $signed(_GEN_11082); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11084 = 10'h34b == cnt[9:0] ? $signed(-32'shd989) : $signed(_GEN_11083); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11085 = 10'h34c == cnt[9:0] ? $signed(-32'shd9f2) : $signed(_GEN_11084); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11086 = 10'h34d == cnt[9:0] ? $signed(-32'shda5c) : $signed(_GEN_11085); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11087 = 10'h34e == cnt[9:0] ? $signed(-32'shdac4) : $signed(_GEN_11086); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11088 = 10'h34f == cnt[9:0] ? $signed(-32'shdb2c) : $signed(_GEN_11087); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11089 = 10'h350 == cnt[9:0] ? $signed(-32'shdb94) : $signed(_GEN_11088); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11090 = 10'h351 == cnt[9:0] ? $signed(-32'shdbfb) : $signed(_GEN_11089); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11091 = 10'h352 == cnt[9:0] ? $signed(-32'shdc62) : $signed(_GEN_11090); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11092 = 10'h353 == cnt[9:0] ? $signed(-32'shdcc8) : $signed(_GEN_11091); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11093 = 10'h354 == cnt[9:0] ? $signed(-32'shdd2d) : $signed(_GEN_11092); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11094 = 10'h355 == cnt[9:0] ? $signed(-32'shdd92) : $signed(_GEN_11093); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11095 = 10'h356 == cnt[9:0] ? $signed(-32'shddf7) : $signed(_GEN_11094); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11096 = 10'h357 == cnt[9:0] ? $signed(-32'shde5b) : $signed(_GEN_11095); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11097 = 10'h358 == cnt[9:0] ? $signed(-32'shdebe) : $signed(_GEN_11096); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11098 = 10'h359 == cnt[9:0] ? $signed(-32'shdf21) : $signed(_GEN_11097); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11099 = 10'h35a == cnt[9:0] ? $signed(-32'shdf83) : $signed(_GEN_11098); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11100 = 10'h35b == cnt[9:0] ? $signed(-32'shdfe5) : $signed(_GEN_11099); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11101 = 10'h35c == cnt[9:0] ? $signed(-32'she046) : $signed(_GEN_11100); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11102 = 10'h35d == cnt[9:0] ? $signed(-32'she0a7) : $signed(_GEN_11101); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11103 = 10'h35e == cnt[9:0] ? $signed(-32'she107) : $signed(_GEN_11102); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11104 = 10'h35f == cnt[9:0] ? $signed(-32'she167) : $signed(_GEN_11103); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11105 = 10'h360 == cnt[9:0] ? $signed(-32'she1c6) : $signed(_GEN_11104); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11106 = 10'h361 == cnt[9:0] ? $signed(-32'she224) : $signed(_GEN_11105); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11107 = 10'h362 == cnt[9:0] ? $signed(-32'she282) : $signed(_GEN_11106); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11108 = 10'h363 == cnt[9:0] ? $signed(-32'she2df) : $signed(_GEN_11107); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11109 = 10'h364 == cnt[9:0] ? $signed(-32'she33c) : $signed(_GEN_11108); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11110 = 10'h365 == cnt[9:0] ? $signed(-32'she399) : $signed(_GEN_11109); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11111 = 10'h366 == cnt[9:0] ? $signed(-32'she3f4) : $signed(_GEN_11110); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11112 = 10'h367 == cnt[9:0] ? $signed(-32'she450) : $signed(_GEN_11111); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11113 = 10'h368 == cnt[9:0] ? $signed(-32'she4aa) : $signed(_GEN_11112); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11114 = 10'h369 == cnt[9:0] ? $signed(-32'she504) : $signed(_GEN_11113); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11115 = 10'h36a == cnt[9:0] ? $signed(-32'she55e) : $signed(_GEN_11114); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11116 = 10'h36b == cnt[9:0] ? $signed(-32'she5b7) : $signed(_GEN_11115); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11117 = 10'h36c == cnt[9:0] ? $signed(-32'she610) : $signed(_GEN_11116); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11118 = 10'h36d == cnt[9:0] ? $signed(-32'she667) : $signed(_GEN_11117); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11119 = 10'h36e == cnt[9:0] ? $signed(-32'she6bf) : $signed(_GEN_11118); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11120 = 10'h36f == cnt[9:0] ? $signed(-32'she716) : $signed(_GEN_11119); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11121 = 10'h370 == cnt[9:0] ? $signed(-32'she76c) : $signed(_GEN_11120); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11122 = 10'h371 == cnt[9:0] ? $signed(-32'she7c2) : $signed(_GEN_11121); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11123 = 10'h372 == cnt[9:0] ? $signed(-32'she817) : $signed(_GEN_11122); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11124 = 10'h373 == cnt[9:0] ? $signed(-32'she86b) : $signed(_GEN_11123); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11125 = 10'h374 == cnt[9:0] ? $signed(-32'she8bf) : $signed(_GEN_11124); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11126 = 10'h375 == cnt[9:0] ? $signed(-32'she913) : $signed(_GEN_11125); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11127 = 10'h376 == cnt[9:0] ? $signed(-32'she966) : $signed(_GEN_11126); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11128 = 10'h377 == cnt[9:0] ? $signed(-32'she9b8) : $signed(_GEN_11127); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11129 = 10'h378 == cnt[9:0] ? $signed(-32'shea0a) : $signed(_GEN_11128); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11130 = 10'h379 == cnt[9:0] ? $signed(-32'shea5b) : $signed(_GEN_11129); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11131 = 10'h37a == cnt[9:0] ? $signed(-32'sheaab) : $signed(_GEN_11130); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11132 = 10'h37b == cnt[9:0] ? $signed(-32'sheafc) : $signed(_GEN_11131); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11133 = 10'h37c == cnt[9:0] ? $signed(-32'sheb4b) : $signed(_GEN_11132); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11134 = 10'h37d == cnt[9:0] ? $signed(-32'sheb9a) : $signed(_GEN_11133); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11135 = 10'h37e == cnt[9:0] ? $signed(-32'shebe8) : $signed(_GEN_11134); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11136 = 10'h37f == cnt[9:0] ? $signed(-32'shec36) : $signed(_GEN_11135); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11137 = 10'h380 == cnt[9:0] ? $signed(-32'shec83) : $signed(_GEN_11136); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11138 = 10'h381 == cnt[9:0] ? $signed(-32'shecd0) : $signed(_GEN_11137); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11139 = 10'h382 == cnt[9:0] ? $signed(-32'shed1c) : $signed(_GEN_11138); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11140 = 10'h383 == cnt[9:0] ? $signed(-32'shed68) : $signed(_GEN_11139); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11141 = 10'h384 == cnt[9:0] ? $signed(-32'shedb3) : $signed(_GEN_11140); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11142 = 10'h385 == cnt[9:0] ? $signed(-32'shedfd) : $signed(_GEN_11141); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11143 = 10'h386 == cnt[9:0] ? $signed(-32'shee47) : $signed(_GEN_11142); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11144 = 10'h387 == cnt[9:0] ? $signed(-32'shee90) : $signed(_GEN_11143); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11145 = 10'h388 == cnt[9:0] ? $signed(-32'sheed9) : $signed(_GEN_11144); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11146 = 10'h389 == cnt[9:0] ? $signed(-32'shef21) : $signed(_GEN_11145); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11147 = 10'h38a == cnt[9:0] ? $signed(-32'shef68) : $signed(_GEN_11146); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11148 = 10'h38b == cnt[9:0] ? $signed(-32'shefaf) : $signed(_GEN_11147); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11149 = 10'h38c == cnt[9:0] ? $signed(-32'sheff5) : $signed(_GEN_11148); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11150 = 10'h38d == cnt[9:0] ? $signed(-32'shf03b) : $signed(_GEN_11149); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11151 = 10'h38e == cnt[9:0] ? $signed(-32'shf080) : $signed(_GEN_11150); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11152 = 10'h38f == cnt[9:0] ? $signed(-32'shf0c5) : $signed(_GEN_11151); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11153 = 10'h390 == cnt[9:0] ? $signed(-32'shf109) : $signed(_GEN_11152); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11154 = 10'h391 == cnt[9:0] ? $signed(-32'shf14c) : $signed(_GEN_11153); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11155 = 10'h392 == cnt[9:0] ? $signed(-32'shf18f) : $signed(_GEN_11154); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11156 = 10'h393 == cnt[9:0] ? $signed(-32'shf1d2) : $signed(_GEN_11155); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11157 = 10'h394 == cnt[9:0] ? $signed(-32'shf213) : $signed(_GEN_11156); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11158 = 10'h395 == cnt[9:0] ? $signed(-32'shf254) : $signed(_GEN_11157); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11159 = 10'h396 == cnt[9:0] ? $signed(-32'shf295) : $signed(_GEN_11158); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11160 = 10'h397 == cnt[9:0] ? $signed(-32'shf2d5) : $signed(_GEN_11159); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11161 = 10'h398 == cnt[9:0] ? $signed(-32'shf314) : $signed(_GEN_11160); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11162 = 10'h399 == cnt[9:0] ? $signed(-32'shf353) : $signed(_GEN_11161); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11163 = 10'h39a == cnt[9:0] ? $signed(-32'shf391) : $signed(_GEN_11162); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11164 = 10'h39b == cnt[9:0] ? $signed(-32'shf3cf) : $signed(_GEN_11163); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11165 = 10'h39c == cnt[9:0] ? $signed(-32'shf40c) : $signed(_GEN_11164); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11166 = 10'h39d == cnt[9:0] ? $signed(-32'shf448) : $signed(_GEN_11165); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11167 = 10'h39e == cnt[9:0] ? $signed(-32'shf484) : $signed(_GEN_11166); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11168 = 10'h39f == cnt[9:0] ? $signed(-32'shf4bf) : $signed(_GEN_11167); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11169 = 10'h3a0 == cnt[9:0] ? $signed(-32'shf4fa) : $signed(_GEN_11168); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11170 = 10'h3a1 == cnt[9:0] ? $signed(-32'shf534) : $signed(_GEN_11169); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11171 = 10'h3a2 == cnt[9:0] ? $signed(-32'shf56e) : $signed(_GEN_11170); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11172 = 10'h3a3 == cnt[9:0] ? $signed(-32'shf5a6) : $signed(_GEN_11171); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11173 = 10'h3a4 == cnt[9:0] ? $signed(-32'shf5df) : $signed(_GEN_11172); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11174 = 10'h3a5 == cnt[9:0] ? $signed(-32'shf616) : $signed(_GEN_11173); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11175 = 10'h3a6 == cnt[9:0] ? $signed(-32'shf64e) : $signed(_GEN_11174); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11176 = 10'h3a7 == cnt[9:0] ? $signed(-32'shf684) : $signed(_GEN_11175); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11177 = 10'h3a8 == cnt[9:0] ? $signed(-32'shf6ba) : $signed(_GEN_11176); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11178 = 10'h3a9 == cnt[9:0] ? $signed(-32'shf6ef) : $signed(_GEN_11177); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11179 = 10'h3aa == cnt[9:0] ? $signed(-32'shf724) : $signed(_GEN_11178); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11180 = 10'h3ab == cnt[9:0] ? $signed(-32'shf758) : $signed(_GEN_11179); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11181 = 10'h3ac == cnt[9:0] ? $signed(-32'shf78c) : $signed(_GEN_11180); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11182 = 10'h3ad == cnt[9:0] ? $signed(-32'shf7bf) : $signed(_GEN_11181); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11183 = 10'h3ae == cnt[9:0] ? $signed(-32'shf7f1) : $signed(_GEN_11182); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11184 = 10'h3af == cnt[9:0] ? $signed(-32'shf823) : $signed(_GEN_11183); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11185 = 10'h3b0 == cnt[9:0] ? $signed(-32'shf854) : $signed(_GEN_11184); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11186 = 10'h3b1 == cnt[9:0] ? $signed(-32'shf885) : $signed(_GEN_11185); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11187 = 10'h3b2 == cnt[9:0] ? $signed(-32'shf8b4) : $signed(_GEN_11186); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11188 = 10'h3b3 == cnt[9:0] ? $signed(-32'shf8e4) : $signed(_GEN_11187); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11189 = 10'h3b4 == cnt[9:0] ? $signed(-32'shf913) : $signed(_GEN_11188); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11190 = 10'h3b5 == cnt[9:0] ? $signed(-32'shf941) : $signed(_GEN_11189); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11191 = 10'h3b6 == cnt[9:0] ? $signed(-32'shf96e) : $signed(_GEN_11190); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11192 = 10'h3b7 == cnt[9:0] ? $signed(-32'shf99b) : $signed(_GEN_11191); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11193 = 10'h3b8 == cnt[9:0] ? $signed(-32'shf9c8) : $signed(_GEN_11192); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11194 = 10'h3b9 == cnt[9:0] ? $signed(-32'shf9f3) : $signed(_GEN_11193); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11195 = 10'h3ba == cnt[9:0] ? $signed(-32'shfa1f) : $signed(_GEN_11194); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11196 = 10'h3bb == cnt[9:0] ? $signed(-32'shfa49) : $signed(_GEN_11195); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11197 = 10'h3bc == cnt[9:0] ? $signed(-32'shfa73) : $signed(_GEN_11196); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11198 = 10'h3bd == cnt[9:0] ? $signed(-32'shfa9c) : $signed(_GEN_11197); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11199 = 10'h3be == cnt[9:0] ? $signed(-32'shfac5) : $signed(_GEN_11198); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11200 = 10'h3bf == cnt[9:0] ? $signed(-32'shfaed) : $signed(_GEN_11199); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11201 = 10'h3c0 == cnt[9:0] ? $signed(-32'shfb15) : $signed(_GEN_11200); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11202 = 10'h3c1 == cnt[9:0] ? $signed(-32'shfb3c) : $signed(_GEN_11201); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11203 = 10'h3c2 == cnt[9:0] ? $signed(-32'shfb62) : $signed(_GEN_11202); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11204 = 10'h3c3 == cnt[9:0] ? $signed(-32'shfb88) : $signed(_GEN_11203); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11205 = 10'h3c4 == cnt[9:0] ? $signed(-32'shfbad) : $signed(_GEN_11204); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11206 = 10'h3c5 == cnt[9:0] ? $signed(-32'shfbd1) : $signed(_GEN_11205); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11207 = 10'h3c6 == cnt[9:0] ? $signed(-32'shfbf5) : $signed(_GEN_11206); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11208 = 10'h3c7 == cnt[9:0] ? $signed(-32'shfc18) : $signed(_GEN_11207); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11209 = 10'h3c8 == cnt[9:0] ? $signed(-32'shfc3b) : $signed(_GEN_11208); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11210 = 10'h3c9 == cnt[9:0] ? $signed(-32'shfc5d) : $signed(_GEN_11209); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11211 = 10'h3ca == cnt[9:0] ? $signed(-32'shfc7f) : $signed(_GEN_11210); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11212 = 10'h3cb == cnt[9:0] ? $signed(-32'shfca0) : $signed(_GEN_11211); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11213 = 10'h3cc == cnt[9:0] ? $signed(-32'shfcc0) : $signed(_GEN_11212); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11214 = 10'h3cd == cnt[9:0] ? $signed(-32'shfcdf) : $signed(_GEN_11213); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11215 = 10'h3ce == cnt[9:0] ? $signed(-32'shfcfe) : $signed(_GEN_11214); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11216 = 10'h3cf == cnt[9:0] ? $signed(-32'shfd1d) : $signed(_GEN_11215); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11217 = 10'h3d0 == cnt[9:0] ? $signed(-32'shfd3b) : $signed(_GEN_11216); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11218 = 10'h3d1 == cnt[9:0] ? $signed(-32'shfd58) : $signed(_GEN_11217); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11219 = 10'h3d2 == cnt[9:0] ? $signed(-32'shfd74) : $signed(_GEN_11218); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11220 = 10'h3d3 == cnt[9:0] ? $signed(-32'shfd90) : $signed(_GEN_11219); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11221 = 10'h3d4 == cnt[9:0] ? $signed(-32'shfdac) : $signed(_GEN_11220); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11222 = 10'h3d5 == cnt[9:0] ? $signed(-32'shfdc7) : $signed(_GEN_11221); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11223 = 10'h3d6 == cnt[9:0] ? $signed(-32'shfde1) : $signed(_GEN_11222); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11224 = 10'h3d7 == cnt[9:0] ? $signed(-32'shfdfa) : $signed(_GEN_11223); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11225 = 10'h3d8 == cnt[9:0] ? $signed(-32'shfe13) : $signed(_GEN_11224); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11226 = 10'h3d9 == cnt[9:0] ? $signed(-32'shfe2b) : $signed(_GEN_11225); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11227 = 10'h3da == cnt[9:0] ? $signed(-32'shfe43) : $signed(_GEN_11226); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11228 = 10'h3db == cnt[9:0] ? $signed(-32'shfe5a) : $signed(_GEN_11227); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11229 = 10'h3dc == cnt[9:0] ? $signed(-32'shfe71) : $signed(_GEN_11228); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11230 = 10'h3dd == cnt[9:0] ? $signed(-32'shfe87) : $signed(_GEN_11229); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11231 = 10'h3de == cnt[9:0] ? $signed(-32'shfe9c) : $signed(_GEN_11230); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11232 = 10'h3df == cnt[9:0] ? $signed(-32'shfeb0) : $signed(_GEN_11231); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11233 = 10'h3e0 == cnt[9:0] ? $signed(-32'shfec4) : $signed(_GEN_11232); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11234 = 10'h3e1 == cnt[9:0] ? $signed(-32'shfed8) : $signed(_GEN_11233); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11235 = 10'h3e2 == cnt[9:0] ? $signed(-32'shfeeb) : $signed(_GEN_11234); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11236 = 10'h3e3 == cnt[9:0] ? $signed(-32'shfefd) : $signed(_GEN_11235); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11237 = 10'h3e4 == cnt[9:0] ? $signed(-32'shff0e) : $signed(_GEN_11236); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11238 = 10'h3e5 == cnt[9:0] ? $signed(-32'shff1f) : $signed(_GEN_11237); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11239 = 10'h3e6 == cnt[9:0] ? $signed(-32'shff30) : $signed(_GEN_11238); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11240 = 10'h3e7 == cnt[9:0] ? $signed(-32'shff3f) : $signed(_GEN_11239); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11241 = 10'h3e8 == cnt[9:0] ? $signed(-32'shff4e) : $signed(_GEN_11240); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11242 = 10'h3e9 == cnt[9:0] ? $signed(-32'shff5d) : $signed(_GEN_11241); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11243 = 10'h3ea == cnt[9:0] ? $signed(-32'shff6b) : $signed(_GEN_11242); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11244 = 10'h3eb == cnt[9:0] ? $signed(-32'shff78) : $signed(_GEN_11243); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11245 = 10'h3ec == cnt[9:0] ? $signed(-32'shff85) : $signed(_GEN_11244); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11246 = 10'h3ed == cnt[9:0] ? $signed(-32'shff91) : $signed(_GEN_11245); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11247 = 10'h3ee == cnt[9:0] ? $signed(-32'shff9c) : $signed(_GEN_11246); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11248 = 10'h3ef == cnt[9:0] ? $signed(-32'shffa7) : $signed(_GEN_11247); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11249 = 10'h3f0 == cnt[9:0] ? $signed(-32'shffb1) : $signed(_GEN_11248); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11250 = 10'h3f1 == cnt[9:0] ? $signed(-32'shffbb) : $signed(_GEN_11249); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11251 = 10'h3f2 == cnt[9:0] ? $signed(-32'shffc4) : $signed(_GEN_11250); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11252 = 10'h3f3 == cnt[9:0] ? $signed(-32'shffcc) : $signed(_GEN_11251); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11253 = 10'h3f4 == cnt[9:0] ? $signed(-32'shffd4) : $signed(_GEN_11252); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11254 = 10'h3f5 == cnt[9:0] ? $signed(-32'shffdb) : $signed(_GEN_11253); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11255 = 10'h3f6 == cnt[9:0] ? $signed(-32'shffe1) : $signed(_GEN_11254); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11256 = 10'h3f7 == cnt[9:0] ? $signed(-32'shffe7) : $signed(_GEN_11255); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11257 = 10'h3f8 == cnt[9:0] ? $signed(-32'shffec) : $signed(_GEN_11256); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11258 = 10'h3f9 == cnt[9:0] ? $signed(-32'shfff1) : $signed(_GEN_11257); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11259 = 10'h3fa == cnt[9:0] ? $signed(-32'shfff5) : $signed(_GEN_11258); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11260 = 10'h3fb == cnt[9:0] ? $signed(-32'shfff8) : $signed(_GEN_11259); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11261 = 10'h3fc == cnt[9:0] ? $signed(-32'shfffb) : $signed(_GEN_11260); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11262 = 10'h3fd == cnt[9:0] ? $signed(-32'shfffd) : $signed(_GEN_11261); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11263 = 10'h3fe == cnt[9:0] ? $signed(-32'shffff) : $signed(_GEN_11262); // @[FFT.scala 34:12]
  wire [31:0] _GEN_11266 = 10'h1 == cnt[9:0] ? $signed(-32'shc9) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11267 = 10'h2 == cnt[9:0] ? $signed(-32'sh192) : $signed(_GEN_11266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11268 = 10'h3 == cnt[9:0] ? $signed(-32'sh25b) : $signed(_GEN_11267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11269 = 10'h4 == cnt[9:0] ? $signed(-32'sh324) : $signed(_GEN_11268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11270 = 10'h5 == cnt[9:0] ? $signed(-32'sh3ed) : $signed(_GEN_11269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11271 = 10'h6 == cnt[9:0] ? $signed(-32'sh4b6) : $signed(_GEN_11270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11272 = 10'h7 == cnt[9:0] ? $signed(-32'sh57f) : $signed(_GEN_11271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11273 = 10'h8 == cnt[9:0] ? $signed(-32'sh648) : $signed(_GEN_11272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11274 = 10'h9 == cnt[9:0] ? $signed(-32'sh711) : $signed(_GEN_11273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11275 = 10'ha == cnt[9:0] ? $signed(-32'sh7da) : $signed(_GEN_11274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11276 = 10'hb == cnt[9:0] ? $signed(-32'sh8a3) : $signed(_GEN_11275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11277 = 10'hc == cnt[9:0] ? $signed(-32'sh96c) : $signed(_GEN_11276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11278 = 10'hd == cnt[9:0] ? $signed(-32'sha35) : $signed(_GEN_11277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11279 = 10'he == cnt[9:0] ? $signed(-32'shafe) : $signed(_GEN_11278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11280 = 10'hf == cnt[9:0] ? $signed(-32'shbc7) : $signed(_GEN_11279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11281 = 10'h10 == cnt[9:0] ? $signed(-32'shc90) : $signed(_GEN_11280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11282 = 10'h11 == cnt[9:0] ? $signed(-32'shd59) : $signed(_GEN_11281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11283 = 10'h12 == cnt[9:0] ? $signed(-32'she21) : $signed(_GEN_11282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11284 = 10'h13 == cnt[9:0] ? $signed(-32'sheea) : $signed(_GEN_11283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11285 = 10'h14 == cnt[9:0] ? $signed(-32'shfb3) : $signed(_GEN_11284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11286 = 10'h15 == cnt[9:0] ? $signed(-32'sh107b) : $signed(_GEN_11285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11287 = 10'h16 == cnt[9:0] ? $signed(-32'sh1144) : $signed(_GEN_11286); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11288 = 10'h17 == cnt[9:0] ? $signed(-32'sh120d) : $signed(_GEN_11287); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11289 = 10'h18 == cnt[9:0] ? $signed(-32'sh12d5) : $signed(_GEN_11288); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11290 = 10'h19 == cnt[9:0] ? $signed(-32'sh139e) : $signed(_GEN_11289); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11291 = 10'h1a == cnt[9:0] ? $signed(-32'sh1466) : $signed(_GEN_11290); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11292 = 10'h1b == cnt[9:0] ? $signed(-32'sh152e) : $signed(_GEN_11291); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11293 = 10'h1c == cnt[9:0] ? $signed(-32'sh15f7) : $signed(_GEN_11292); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11294 = 10'h1d == cnt[9:0] ? $signed(-32'sh16bf) : $signed(_GEN_11293); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11295 = 10'h1e == cnt[9:0] ? $signed(-32'sh1787) : $signed(_GEN_11294); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11296 = 10'h1f == cnt[9:0] ? $signed(-32'sh1850) : $signed(_GEN_11295); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11297 = 10'h20 == cnt[9:0] ? $signed(-32'sh1918) : $signed(_GEN_11296); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11298 = 10'h21 == cnt[9:0] ? $signed(-32'sh19e0) : $signed(_GEN_11297); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11299 = 10'h22 == cnt[9:0] ? $signed(-32'sh1aa8) : $signed(_GEN_11298); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11300 = 10'h23 == cnt[9:0] ? $signed(-32'sh1b70) : $signed(_GEN_11299); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11301 = 10'h24 == cnt[9:0] ? $signed(-32'sh1c38) : $signed(_GEN_11300); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11302 = 10'h25 == cnt[9:0] ? $signed(-32'sh1cff) : $signed(_GEN_11301); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11303 = 10'h26 == cnt[9:0] ? $signed(-32'sh1dc7) : $signed(_GEN_11302); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11304 = 10'h27 == cnt[9:0] ? $signed(-32'sh1e8f) : $signed(_GEN_11303); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11305 = 10'h28 == cnt[9:0] ? $signed(-32'sh1f56) : $signed(_GEN_11304); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11306 = 10'h29 == cnt[9:0] ? $signed(-32'sh201e) : $signed(_GEN_11305); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11307 = 10'h2a == cnt[9:0] ? $signed(-32'sh20e5) : $signed(_GEN_11306); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11308 = 10'h2b == cnt[9:0] ? $signed(-32'sh21ad) : $signed(_GEN_11307); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11309 = 10'h2c == cnt[9:0] ? $signed(-32'sh2274) : $signed(_GEN_11308); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11310 = 10'h2d == cnt[9:0] ? $signed(-32'sh233b) : $signed(_GEN_11309); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11311 = 10'h2e == cnt[9:0] ? $signed(-32'sh2402) : $signed(_GEN_11310); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11312 = 10'h2f == cnt[9:0] ? $signed(-32'sh24c9) : $signed(_GEN_11311); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11313 = 10'h30 == cnt[9:0] ? $signed(-32'sh2590) : $signed(_GEN_11312); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11314 = 10'h31 == cnt[9:0] ? $signed(-32'sh2657) : $signed(_GEN_11313); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11315 = 10'h32 == cnt[9:0] ? $signed(-32'sh271e) : $signed(_GEN_11314); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11316 = 10'h33 == cnt[9:0] ? $signed(-32'sh27e4) : $signed(_GEN_11315); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11317 = 10'h34 == cnt[9:0] ? $signed(-32'sh28ab) : $signed(_GEN_11316); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11318 = 10'h35 == cnt[9:0] ? $signed(-32'sh2971) : $signed(_GEN_11317); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11319 = 10'h36 == cnt[9:0] ? $signed(-32'sh2a38) : $signed(_GEN_11318); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11320 = 10'h37 == cnt[9:0] ? $signed(-32'sh2afe) : $signed(_GEN_11319); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11321 = 10'h38 == cnt[9:0] ? $signed(-32'sh2bc4) : $signed(_GEN_11320); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11322 = 10'h39 == cnt[9:0] ? $signed(-32'sh2c8a) : $signed(_GEN_11321); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11323 = 10'h3a == cnt[9:0] ? $signed(-32'sh2d50) : $signed(_GEN_11322); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11324 = 10'h3b == cnt[9:0] ? $signed(-32'sh2e16) : $signed(_GEN_11323); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11325 = 10'h3c == cnt[9:0] ? $signed(-32'sh2edc) : $signed(_GEN_11324); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11326 = 10'h3d == cnt[9:0] ? $signed(-32'sh2fa1) : $signed(_GEN_11325); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11327 = 10'h3e == cnt[9:0] ? $signed(-32'sh3067) : $signed(_GEN_11326); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11328 = 10'h3f == cnt[9:0] ? $signed(-32'sh312c) : $signed(_GEN_11327); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11329 = 10'h40 == cnt[9:0] ? $signed(-32'sh31f1) : $signed(_GEN_11328); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11330 = 10'h41 == cnt[9:0] ? $signed(-32'sh32b7) : $signed(_GEN_11329); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11331 = 10'h42 == cnt[9:0] ? $signed(-32'sh337c) : $signed(_GEN_11330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11332 = 10'h43 == cnt[9:0] ? $signed(-32'sh3440) : $signed(_GEN_11331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11333 = 10'h44 == cnt[9:0] ? $signed(-32'sh3505) : $signed(_GEN_11332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11334 = 10'h45 == cnt[9:0] ? $signed(-32'sh35ca) : $signed(_GEN_11333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11335 = 10'h46 == cnt[9:0] ? $signed(-32'sh368e) : $signed(_GEN_11334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11336 = 10'h47 == cnt[9:0] ? $signed(-32'sh3753) : $signed(_GEN_11335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11337 = 10'h48 == cnt[9:0] ? $signed(-32'sh3817) : $signed(_GEN_11336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11338 = 10'h49 == cnt[9:0] ? $signed(-32'sh38db) : $signed(_GEN_11337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11339 = 10'h4a == cnt[9:0] ? $signed(-32'sh399f) : $signed(_GEN_11338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11340 = 10'h4b == cnt[9:0] ? $signed(-32'sh3a63) : $signed(_GEN_11339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11341 = 10'h4c == cnt[9:0] ? $signed(-32'sh3b27) : $signed(_GEN_11340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11342 = 10'h4d == cnt[9:0] ? $signed(-32'sh3bea) : $signed(_GEN_11341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11343 = 10'h4e == cnt[9:0] ? $signed(-32'sh3cae) : $signed(_GEN_11342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11344 = 10'h4f == cnt[9:0] ? $signed(-32'sh3d71) : $signed(_GEN_11343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11345 = 10'h50 == cnt[9:0] ? $signed(-32'sh3e34) : $signed(_GEN_11344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11346 = 10'h51 == cnt[9:0] ? $signed(-32'sh3ef7) : $signed(_GEN_11345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11347 = 10'h52 == cnt[9:0] ? $signed(-32'sh3fba) : $signed(_GEN_11346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11348 = 10'h53 == cnt[9:0] ? $signed(-32'sh407c) : $signed(_GEN_11347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11349 = 10'h54 == cnt[9:0] ? $signed(-32'sh413f) : $signed(_GEN_11348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11350 = 10'h55 == cnt[9:0] ? $signed(-32'sh4201) : $signed(_GEN_11349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11351 = 10'h56 == cnt[9:0] ? $signed(-32'sh42c3) : $signed(_GEN_11350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11352 = 10'h57 == cnt[9:0] ? $signed(-32'sh4385) : $signed(_GEN_11351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11353 = 10'h58 == cnt[9:0] ? $signed(-32'sh4447) : $signed(_GEN_11352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11354 = 10'h59 == cnt[9:0] ? $signed(-32'sh4509) : $signed(_GEN_11353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11355 = 10'h5a == cnt[9:0] ? $signed(-32'sh45cb) : $signed(_GEN_11354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11356 = 10'h5b == cnt[9:0] ? $signed(-32'sh468c) : $signed(_GEN_11355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11357 = 10'h5c == cnt[9:0] ? $signed(-32'sh474d) : $signed(_GEN_11356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11358 = 10'h5d == cnt[9:0] ? $signed(-32'sh480e) : $signed(_GEN_11357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11359 = 10'h5e == cnt[9:0] ? $signed(-32'sh48cf) : $signed(_GEN_11358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11360 = 10'h5f == cnt[9:0] ? $signed(-32'sh4990) : $signed(_GEN_11359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11361 = 10'h60 == cnt[9:0] ? $signed(-32'sh4a50) : $signed(_GEN_11360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11362 = 10'h61 == cnt[9:0] ? $signed(-32'sh4b10) : $signed(_GEN_11361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11363 = 10'h62 == cnt[9:0] ? $signed(-32'sh4bd1) : $signed(_GEN_11362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11364 = 10'h63 == cnt[9:0] ? $signed(-32'sh4c90) : $signed(_GEN_11363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11365 = 10'h64 == cnt[9:0] ? $signed(-32'sh4d50) : $signed(_GEN_11364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11366 = 10'h65 == cnt[9:0] ? $signed(-32'sh4e10) : $signed(_GEN_11365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11367 = 10'h66 == cnt[9:0] ? $signed(-32'sh4ecf) : $signed(_GEN_11366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11368 = 10'h67 == cnt[9:0] ? $signed(-32'sh4f8e) : $signed(_GEN_11367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11369 = 10'h68 == cnt[9:0] ? $signed(-32'sh504d) : $signed(_GEN_11368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11370 = 10'h69 == cnt[9:0] ? $signed(-32'sh510c) : $signed(_GEN_11369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11371 = 10'h6a == cnt[9:0] ? $signed(-32'sh51cb) : $signed(_GEN_11370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11372 = 10'h6b == cnt[9:0] ? $signed(-32'sh5289) : $signed(_GEN_11371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11373 = 10'h6c == cnt[9:0] ? $signed(-32'sh5348) : $signed(_GEN_11372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11374 = 10'h6d == cnt[9:0] ? $signed(-32'sh5406) : $signed(_GEN_11373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11375 = 10'h6e == cnt[9:0] ? $signed(-32'sh54c3) : $signed(_GEN_11374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11376 = 10'h6f == cnt[9:0] ? $signed(-32'sh5581) : $signed(_GEN_11375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11377 = 10'h70 == cnt[9:0] ? $signed(-32'sh563e) : $signed(_GEN_11376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11378 = 10'h71 == cnt[9:0] ? $signed(-32'sh56fc) : $signed(_GEN_11377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11379 = 10'h72 == cnt[9:0] ? $signed(-32'sh57b9) : $signed(_GEN_11378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11380 = 10'h73 == cnt[9:0] ? $signed(-32'sh5875) : $signed(_GEN_11379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11381 = 10'h74 == cnt[9:0] ? $signed(-32'sh5932) : $signed(_GEN_11380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11382 = 10'h75 == cnt[9:0] ? $signed(-32'sh59ee) : $signed(_GEN_11381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11383 = 10'h76 == cnt[9:0] ? $signed(-32'sh5aaa) : $signed(_GEN_11382); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11384 = 10'h77 == cnt[9:0] ? $signed(-32'sh5b66) : $signed(_GEN_11383); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11385 = 10'h78 == cnt[9:0] ? $signed(-32'sh5c22) : $signed(_GEN_11384); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11386 = 10'h79 == cnt[9:0] ? $signed(-32'sh5cde) : $signed(_GEN_11385); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11387 = 10'h7a == cnt[9:0] ? $signed(-32'sh5d99) : $signed(_GEN_11386); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11388 = 10'h7b == cnt[9:0] ? $signed(-32'sh5e54) : $signed(_GEN_11387); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11389 = 10'h7c == cnt[9:0] ? $signed(-32'sh5f0f) : $signed(_GEN_11388); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11390 = 10'h7d == cnt[9:0] ? $signed(-32'sh5fc9) : $signed(_GEN_11389); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11391 = 10'h7e == cnt[9:0] ? $signed(-32'sh6084) : $signed(_GEN_11390); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11392 = 10'h7f == cnt[9:0] ? $signed(-32'sh613e) : $signed(_GEN_11391); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11393 = 10'h80 == cnt[9:0] ? $signed(-32'sh61f8) : $signed(_GEN_11392); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11394 = 10'h81 == cnt[9:0] ? $signed(-32'sh62b1) : $signed(_GEN_11393); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11395 = 10'h82 == cnt[9:0] ? $signed(-32'sh636b) : $signed(_GEN_11394); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11396 = 10'h83 == cnt[9:0] ? $signed(-32'sh6424) : $signed(_GEN_11395); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11397 = 10'h84 == cnt[9:0] ? $signed(-32'sh64dd) : $signed(_GEN_11396); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11398 = 10'h85 == cnt[9:0] ? $signed(-32'sh6595) : $signed(_GEN_11397); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11399 = 10'h86 == cnt[9:0] ? $signed(-32'sh664e) : $signed(_GEN_11398); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11400 = 10'h87 == cnt[9:0] ? $signed(-32'sh6706) : $signed(_GEN_11399); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11401 = 10'h88 == cnt[9:0] ? $signed(-32'sh67be) : $signed(_GEN_11400); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11402 = 10'h89 == cnt[9:0] ? $signed(-32'sh6876) : $signed(_GEN_11401); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11403 = 10'h8a == cnt[9:0] ? $signed(-32'sh692d) : $signed(_GEN_11402); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11404 = 10'h8b == cnt[9:0] ? $signed(-32'sh69e4) : $signed(_GEN_11403); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11405 = 10'h8c == cnt[9:0] ? $signed(-32'sh6a9b) : $signed(_GEN_11404); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11406 = 10'h8d == cnt[9:0] ? $signed(-32'sh6b52) : $signed(_GEN_11405); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11407 = 10'h8e == cnt[9:0] ? $signed(-32'sh6c08) : $signed(_GEN_11406); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11408 = 10'h8f == cnt[9:0] ? $signed(-32'sh6cbe) : $signed(_GEN_11407); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11409 = 10'h90 == cnt[9:0] ? $signed(-32'sh6d74) : $signed(_GEN_11408); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11410 = 10'h91 == cnt[9:0] ? $signed(-32'sh6e2a) : $signed(_GEN_11409); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11411 = 10'h92 == cnt[9:0] ? $signed(-32'sh6edf) : $signed(_GEN_11410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11412 = 10'h93 == cnt[9:0] ? $signed(-32'sh6f94) : $signed(_GEN_11411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11413 = 10'h94 == cnt[9:0] ? $signed(-32'sh7049) : $signed(_GEN_11412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11414 = 10'h95 == cnt[9:0] ? $signed(-32'sh70fe) : $signed(_GEN_11413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11415 = 10'h96 == cnt[9:0] ? $signed(-32'sh71b2) : $signed(_GEN_11414); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11416 = 10'h97 == cnt[9:0] ? $signed(-32'sh7266) : $signed(_GEN_11415); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11417 = 10'h98 == cnt[9:0] ? $signed(-32'sh731a) : $signed(_GEN_11416); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11418 = 10'h99 == cnt[9:0] ? $signed(-32'sh73cd) : $signed(_GEN_11417); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11419 = 10'h9a == cnt[9:0] ? $signed(-32'sh7480) : $signed(_GEN_11418); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11420 = 10'h9b == cnt[9:0] ? $signed(-32'sh7533) : $signed(_GEN_11419); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11421 = 10'h9c == cnt[9:0] ? $signed(-32'sh75e6) : $signed(_GEN_11420); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11422 = 10'h9d == cnt[9:0] ? $signed(-32'sh7698) : $signed(_GEN_11421); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11423 = 10'h9e == cnt[9:0] ? $signed(-32'sh774a) : $signed(_GEN_11422); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11424 = 10'h9f == cnt[9:0] ? $signed(-32'sh77fc) : $signed(_GEN_11423); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11425 = 10'ha0 == cnt[9:0] ? $signed(-32'sh78ad) : $signed(_GEN_11424); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11426 = 10'ha1 == cnt[9:0] ? $signed(-32'sh795f) : $signed(_GEN_11425); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11427 = 10'ha2 == cnt[9:0] ? $signed(-32'sh7a10) : $signed(_GEN_11426); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11428 = 10'ha3 == cnt[9:0] ? $signed(-32'sh7ac0) : $signed(_GEN_11427); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11429 = 10'ha4 == cnt[9:0] ? $signed(-32'sh7b70) : $signed(_GEN_11428); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11430 = 10'ha5 == cnt[9:0] ? $signed(-32'sh7c20) : $signed(_GEN_11429); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11431 = 10'ha6 == cnt[9:0] ? $signed(-32'sh7cd0) : $signed(_GEN_11430); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11432 = 10'ha7 == cnt[9:0] ? $signed(-32'sh7d7f) : $signed(_GEN_11431); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11433 = 10'ha8 == cnt[9:0] ? $signed(-32'sh7e2f) : $signed(_GEN_11432); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11434 = 10'ha9 == cnt[9:0] ? $signed(-32'sh7edd) : $signed(_GEN_11433); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11435 = 10'haa == cnt[9:0] ? $signed(-32'sh7f8c) : $signed(_GEN_11434); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11436 = 10'hab == cnt[9:0] ? $signed(-32'sh803a) : $signed(_GEN_11435); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11437 = 10'hac == cnt[9:0] ? $signed(-32'sh80e8) : $signed(_GEN_11436); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11438 = 10'had == cnt[9:0] ? $signed(-32'sh8195) : $signed(_GEN_11437); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11439 = 10'hae == cnt[9:0] ? $signed(-32'sh8243) : $signed(_GEN_11438); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11440 = 10'haf == cnt[9:0] ? $signed(-32'sh82f0) : $signed(_GEN_11439); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11441 = 10'hb0 == cnt[9:0] ? $signed(-32'sh839c) : $signed(_GEN_11440); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11442 = 10'hb1 == cnt[9:0] ? $signed(-32'sh8449) : $signed(_GEN_11441); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11443 = 10'hb2 == cnt[9:0] ? $signed(-32'sh84f5) : $signed(_GEN_11442); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11444 = 10'hb3 == cnt[9:0] ? $signed(-32'sh85a0) : $signed(_GEN_11443); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11445 = 10'hb4 == cnt[9:0] ? $signed(-32'sh864c) : $signed(_GEN_11444); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11446 = 10'hb5 == cnt[9:0] ? $signed(-32'sh86f7) : $signed(_GEN_11445); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11447 = 10'hb6 == cnt[9:0] ? $signed(-32'sh87a1) : $signed(_GEN_11446); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11448 = 10'hb7 == cnt[9:0] ? $signed(-32'sh884c) : $signed(_GEN_11447); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11449 = 10'hb8 == cnt[9:0] ? $signed(-32'sh88f6) : $signed(_GEN_11448); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11450 = 10'hb9 == cnt[9:0] ? $signed(-32'sh899f) : $signed(_GEN_11449); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11451 = 10'hba == cnt[9:0] ? $signed(-32'sh8a49) : $signed(_GEN_11450); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11452 = 10'hbb == cnt[9:0] ? $signed(-32'sh8af2) : $signed(_GEN_11451); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11453 = 10'hbc == cnt[9:0] ? $signed(-32'sh8b9a) : $signed(_GEN_11452); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11454 = 10'hbd == cnt[9:0] ? $signed(-32'sh8c43) : $signed(_GEN_11453); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11455 = 10'hbe == cnt[9:0] ? $signed(-32'sh8ceb) : $signed(_GEN_11454); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11456 = 10'hbf == cnt[9:0] ? $signed(-32'sh8d93) : $signed(_GEN_11455); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11457 = 10'hc0 == cnt[9:0] ? $signed(-32'sh8e3a) : $signed(_GEN_11456); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11458 = 10'hc1 == cnt[9:0] ? $signed(-32'sh8ee1) : $signed(_GEN_11457); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11459 = 10'hc2 == cnt[9:0] ? $signed(-32'sh8f88) : $signed(_GEN_11458); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11460 = 10'hc3 == cnt[9:0] ? $signed(-32'sh902e) : $signed(_GEN_11459); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11461 = 10'hc4 == cnt[9:0] ? $signed(-32'sh90d4) : $signed(_GEN_11460); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11462 = 10'hc5 == cnt[9:0] ? $signed(-32'sh9179) : $signed(_GEN_11461); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11463 = 10'hc6 == cnt[9:0] ? $signed(-32'sh921f) : $signed(_GEN_11462); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11464 = 10'hc7 == cnt[9:0] ? $signed(-32'sh92c4) : $signed(_GEN_11463); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11465 = 10'hc8 == cnt[9:0] ? $signed(-32'sh9368) : $signed(_GEN_11464); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11466 = 10'hc9 == cnt[9:0] ? $signed(-32'sh940c) : $signed(_GEN_11465); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11467 = 10'hca == cnt[9:0] ? $signed(-32'sh94b0) : $signed(_GEN_11466); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11468 = 10'hcb == cnt[9:0] ? $signed(-32'sh9554) : $signed(_GEN_11467); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11469 = 10'hcc == cnt[9:0] ? $signed(-32'sh95f7) : $signed(_GEN_11468); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11470 = 10'hcd == cnt[9:0] ? $signed(-32'sh969a) : $signed(_GEN_11469); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11471 = 10'hce == cnt[9:0] ? $signed(-32'sh973c) : $signed(_GEN_11470); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11472 = 10'hcf == cnt[9:0] ? $signed(-32'sh97de) : $signed(_GEN_11471); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11473 = 10'hd0 == cnt[9:0] ? $signed(-32'sh9880) : $signed(_GEN_11472); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11474 = 10'hd1 == cnt[9:0] ? $signed(-32'sh9921) : $signed(_GEN_11473); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11475 = 10'hd2 == cnt[9:0] ? $signed(-32'sh99c2) : $signed(_GEN_11474); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11476 = 10'hd3 == cnt[9:0] ? $signed(-32'sh9a63) : $signed(_GEN_11475); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11477 = 10'hd4 == cnt[9:0] ? $signed(-32'sh9b03) : $signed(_GEN_11476); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11478 = 10'hd5 == cnt[9:0] ? $signed(-32'sh9ba3) : $signed(_GEN_11477); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11479 = 10'hd6 == cnt[9:0] ? $signed(-32'sh9c42) : $signed(_GEN_11478); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11480 = 10'hd7 == cnt[9:0] ? $signed(-32'sh9ce1) : $signed(_GEN_11479); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11481 = 10'hd8 == cnt[9:0] ? $signed(-32'sh9d80) : $signed(_GEN_11480); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11482 = 10'hd9 == cnt[9:0] ? $signed(-32'sh9e1e) : $signed(_GEN_11481); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11483 = 10'hda == cnt[9:0] ? $signed(-32'sh9ebc) : $signed(_GEN_11482); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11484 = 10'hdb == cnt[9:0] ? $signed(-32'sh9f5a) : $signed(_GEN_11483); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11485 = 10'hdc == cnt[9:0] ? $signed(-32'sh9ff7) : $signed(_GEN_11484); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11486 = 10'hdd == cnt[9:0] ? $signed(-32'sha094) : $signed(_GEN_11485); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11487 = 10'hde == cnt[9:0] ? $signed(-32'sha130) : $signed(_GEN_11486); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11488 = 10'hdf == cnt[9:0] ? $signed(-32'sha1cc) : $signed(_GEN_11487); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11489 = 10'he0 == cnt[9:0] ? $signed(-32'sha268) : $signed(_GEN_11488); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11490 = 10'he1 == cnt[9:0] ? $signed(-32'sha303) : $signed(_GEN_11489); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11491 = 10'he2 == cnt[9:0] ? $signed(-32'sha39e) : $signed(_GEN_11490); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11492 = 10'he3 == cnt[9:0] ? $signed(-32'sha438) : $signed(_GEN_11491); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11493 = 10'he4 == cnt[9:0] ? $signed(-32'sha4d2) : $signed(_GEN_11492); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11494 = 10'he5 == cnt[9:0] ? $signed(-32'sha56c) : $signed(_GEN_11493); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11495 = 10'he6 == cnt[9:0] ? $signed(-32'sha605) : $signed(_GEN_11494); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11496 = 10'he7 == cnt[9:0] ? $signed(-32'sha69e) : $signed(_GEN_11495); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11497 = 10'he8 == cnt[9:0] ? $signed(-32'sha736) : $signed(_GEN_11496); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11498 = 10'he9 == cnt[9:0] ? $signed(-32'sha7ce) : $signed(_GEN_11497); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11499 = 10'hea == cnt[9:0] ? $signed(-32'sha866) : $signed(_GEN_11498); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11500 = 10'heb == cnt[9:0] ? $signed(-32'sha8fd) : $signed(_GEN_11499); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11501 = 10'hec == cnt[9:0] ? $signed(-32'sha994) : $signed(_GEN_11500); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11502 = 10'hed == cnt[9:0] ? $signed(-32'shaa2a) : $signed(_GEN_11501); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11503 = 10'hee == cnt[9:0] ? $signed(-32'shaac1) : $signed(_GEN_11502); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11504 = 10'hef == cnt[9:0] ? $signed(-32'shab56) : $signed(_GEN_11503); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11505 = 10'hf0 == cnt[9:0] ? $signed(-32'shabeb) : $signed(_GEN_11504); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11506 = 10'hf1 == cnt[9:0] ? $signed(-32'shac80) : $signed(_GEN_11505); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11507 = 10'hf2 == cnt[9:0] ? $signed(-32'shad14) : $signed(_GEN_11506); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11508 = 10'hf3 == cnt[9:0] ? $signed(-32'shada8) : $signed(_GEN_11507); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11509 = 10'hf4 == cnt[9:0] ? $signed(-32'shae3c) : $signed(_GEN_11508); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11510 = 10'hf5 == cnt[9:0] ? $signed(-32'shaecf) : $signed(_GEN_11509); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11511 = 10'hf6 == cnt[9:0] ? $signed(-32'shaf62) : $signed(_GEN_11510); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11512 = 10'hf7 == cnt[9:0] ? $signed(-32'shaff4) : $signed(_GEN_11511); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11513 = 10'hf8 == cnt[9:0] ? $signed(-32'shb086) : $signed(_GEN_11512); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11514 = 10'hf9 == cnt[9:0] ? $signed(-32'shb117) : $signed(_GEN_11513); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11515 = 10'hfa == cnt[9:0] ? $signed(-32'shb1a8) : $signed(_GEN_11514); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11516 = 10'hfb == cnt[9:0] ? $signed(-32'shb239) : $signed(_GEN_11515); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11517 = 10'hfc == cnt[9:0] ? $signed(-32'shb2c9) : $signed(_GEN_11516); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11518 = 10'hfd == cnt[9:0] ? $signed(-32'shb358) : $signed(_GEN_11517); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11519 = 10'hfe == cnt[9:0] ? $signed(-32'shb3e8) : $signed(_GEN_11518); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11520 = 10'hff == cnt[9:0] ? $signed(-32'shb477) : $signed(_GEN_11519); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11521 = 10'h100 == cnt[9:0] ? $signed(-32'shb505) : $signed(_GEN_11520); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11522 = 10'h101 == cnt[9:0] ? $signed(-32'shb593) : $signed(_GEN_11521); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11523 = 10'h102 == cnt[9:0] ? $signed(-32'shb620) : $signed(_GEN_11522); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11524 = 10'h103 == cnt[9:0] ? $signed(-32'shb6ad) : $signed(_GEN_11523); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11525 = 10'h104 == cnt[9:0] ? $signed(-32'shb73a) : $signed(_GEN_11524); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11526 = 10'h105 == cnt[9:0] ? $signed(-32'shb7c6) : $signed(_GEN_11525); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11527 = 10'h106 == cnt[9:0] ? $signed(-32'shb852) : $signed(_GEN_11526); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11528 = 10'h107 == cnt[9:0] ? $signed(-32'shb8dd) : $signed(_GEN_11527); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11529 = 10'h108 == cnt[9:0] ? $signed(-32'shb968) : $signed(_GEN_11528); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11530 = 10'h109 == cnt[9:0] ? $signed(-32'shb9f3) : $signed(_GEN_11529); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11531 = 10'h10a == cnt[9:0] ? $signed(-32'shba7d) : $signed(_GEN_11530); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11532 = 10'h10b == cnt[9:0] ? $signed(-32'shbb06) : $signed(_GEN_11531); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11533 = 10'h10c == cnt[9:0] ? $signed(-32'shbb8f) : $signed(_GEN_11532); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11534 = 10'h10d == cnt[9:0] ? $signed(-32'shbc18) : $signed(_GEN_11533); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11535 = 10'h10e == cnt[9:0] ? $signed(-32'shbca0) : $signed(_GEN_11534); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11536 = 10'h10f == cnt[9:0] ? $signed(-32'shbd28) : $signed(_GEN_11535); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11537 = 10'h110 == cnt[9:0] ? $signed(-32'shbdaf) : $signed(_GEN_11536); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11538 = 10'h111 == cnt[9:0] ? $signed(-32'shbe36) : $signed(_GEN_11537); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11539 = 10'h112 == cnt[9:0] ? $signed(-32'shbebc) : $signed(_GEN_11538); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11540 = 10'h113 == cnt[9:0] ? $signed(-32'shbf42) : $signed(_GEN_11539); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11541 = 10'h114 == cnt[9:0] ? $signed(-32'shbfc7) : $signed(_GEN_11540); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11542 = 10'h115 == cnt[9:0] ? $signed(-32'shc04c) : $signed(_GEN_11541); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11543 = 10'h116 == cnt[9:0] ? $signed(-32'shc0d1) : $signed(_GEN_11542); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11544 = 10'h117 == cnt[9:0] ? $signed(-32'shc155) : $signed(_GEN_11543); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11545 = 10'h118 == cnt[9:0] ? $signed(-32'shc1d8) : $signed(_GEN_11544); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11546 = 10'h119 == cnt[9:0] ? $signed(-32'shc25c) : $signed(_GEN_11545); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11547 = 10'h11a == cnt[9:0] ? $signed(-32'shc2de) : $signed(_GEN_11546); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11548 = 10'h11b == cnt[9:0] ? $signed(-32'shc360) : $signed(_GEN_11547); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11549 = 10'h11c == cnt[9:0] ? $signed(-32'shc3e2) : $signed(_GEN_11548); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11550 = 10'h11d == cnt[9:0] ? $signed(-32'shc463) : $signed(_GEN_11549); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11551 = 10'h11e == cnt[9:0] ? $signed(-32'shc4e4) : $signed(_GEN_11550); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11552 = 10'h11f == cnt[9:0] ? $signed(-32'shc564) : $signed(_GEN_11551); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11553 = 10'h120 == cnt[9:0] ? $signed(-32'shc5e4) : $signed(_GEN_11552); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11554 = 10'h121 == cnt[9:0] ? $signed(-32'shc663) : $signed(_GEN_11553); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11555 = 10'h122 == cnt[9:0] ? $signed(-32'shc6e2) : $signed(_GEN_11554); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11556 = 10'h123 == cnt[9:0] ? $signed(-32'shc761) : $signed(_GEN_11555); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11557 = 10'h124 == cnt[9:0] ? $signed(-32'shc7de) : $signed(_GEN_11556); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11558 = 10'h125 == cnt[9:0] ? $signed(-32'shc85c) : $signed(_GEN_11557); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11559 = 10'h126 == cnt[9:0] ? $signed(-32'shc8d9) : $signed(_GEN_11558); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11560 = 10'h127 == cnt[9:0] ? $signed(-32'shc955) : $signed(_GEN_11559); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11561 = 10'h128 == cnt[9:0] ? $signed(-32'shc9d1) : $signed(_GEN_11560); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11562 = 10'h129 == cnt[9:0] ? $signed(-32'shca4d) : $signed(_GEN_11561); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11563 = 10'h12a == cnt[9:0] ? $signed(-32'shcac7) : $signed(_GEN_11562); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11564 = 10'h12b == cnt[9:0] ? $signed(-32'shcb42) : $signed(_GEN_11563); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11565 = 10'h12c == cnt[9:0] ? $signed(-32'shcbbc) : $signed(_GEN_11564); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11566 = 10'h12d == cnt[9:0] ? $signed(-32'shcc35) : $signed(_GEN_11565); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11567 = 10'h12e == cnt[9:0] ? $signed(-32'shccae) : $signed(_GEN_11566); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11568 = 10'h12f == cnt[9:0] ? $signed(-32'shcd27) : $signed(_GEN_11567); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11569 = 10'h130 == cnt[9:0] ? $signed(-32'shcd9f) : $signed(_GEN_11568); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11570 = 10'h131 == cnt[9:0] ? $signed(-32'shce17) : $signed(_GEN_11569); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11571 = 10'h132 == cnt[9:0] ? $signed(-32'shce8e) : $signed(_GEN_11570); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11572 = 10'h133 == cnt[9:0] ? $signed(-32'shcf04) : $signed(_GEN_11571); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11573 = 10'h134 == cnt[9:0] ? $signed(-32'shcf7a) : $signed(_GEN_11572); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11574 = 10'h135 == cnt[9:0] ? $signed(-32'shcff0) : $signed(_GEN_11573); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11575 = 10'h136 == cnt[9:0] ? $signed(-32'shd065) : $signed(_GEN_11574); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11576 = 10'h137 == cnt[9:0] ? $signed(-32'shd0d9) : $signed(_GEN_11575); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11577 = 10'h138 == cnt[9:0] ? $signed(-32'shd14d) : $signed(_GEN_11576); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11578 = 10'h139 == cnt[9:0] ? $signed(-32'shd1c1) : $signed(_GEN_11577); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11579 = 10'h13a == cnt[9:0] ? $signed(-32'shd234) : $signed(_GEN_11578); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11580 = 10'h13b == cnt[9:0] ? $signed(-32'shd2a6) : $signed(_GEN_11579); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11581 = 10'h13c == cnt[9:0] ? $signed(-32'shd318) : $signed(_GEN_11580); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11582 = 10'h13d == cnt[9:0] ? $signed(-32'shd38a) : $signed(_GEN_11581); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11583 = 10'h13e == cnt[9:0] ? $signed(-32'shd3fb) : $signed(_GEN_11582); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11584 = 10'h13f == cnt[9:0] ? $signed(-32'shd46b) : $signed(_GEN_11583); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11585 = 10'h140 == cnt[9:0] ? $signed(-32'shd4db) : $signed(_GEN_11584); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11586 = 10'h141 == cnt[9:0] ? $signed(-32'shd54b) : $signed(_GEN_11585); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11587 = 10'h142 == cnt[9:0] ? $signed(-32'shd5ba) : $signed(_GEN_11586); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11588 = 10'h143 == cnt[9:0] ? $signed(-32'shd628) : $signed(_GEN_11587); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11589 = 10'h144 == cnt[9:0] ? $signed(-32'shd696) : $signed(_GEN_11588); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11590 = 10'h145 == cnt[9:0] ? $signed(-32'shd703) : $signed(_GEN_11589); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11591 = 10'h146 == cnt[9:0] ? $signed(-32'shd770) : $signed(_GEN_11590); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11592 = 10'h147 == cnt[9:0] ? $signed(-32'shd7dc) : $signed(_GEN_11591); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11593 = 10'h148 == cnt[9:0] ? $signed(-32'shd848) : $signed(_GEN_11592); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11594 = 10'h149 == cnt[9:0] ? $signed(-32'shd8b4) : $signed(_GEN_11593); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11595 = 10'h14a == cnt[9:0] ? $signed(-32'shd91e) : $signed(_GEN_11594); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11596 = 10'h14b == cnt[9:0] ? $signed(-32'shd989) : $signed(_GEN_11595); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11597 = 10'h14c == cnt[9:0] ? $signed(-32'shd9f2) : $signed(_GEN_11596); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11598 = 10'h14d == cnt[9:0] ? $signed(-32'shda5c) : $signed(_GEN_11597); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11599 = 10'h14e == cnt[9:0] ? $signed(-32'shdac4) : $signed(_GEN_11598); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11600 = 10'h14f == cnt[9:0] ? $signed(-32'shdb2c) : $signed(_GEN_11599); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11601 = 10'h150 == cnt[9:0] ? $signed(-32'shdb94) : $signed(_GEN_11600); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11602 = 10'h151 == cnt[9:0] ? $signed(-32'shdbfb) : $signed(_GEN_11601); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11603 = 10'h152 == cnt[9:0] ? $signed(-32'shdc62) : $signed(_GEN_11602); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11604 = 10'h153 == cnt[9:0] ? $signed(-32'shdcc8) : $signed(_GEN_11603); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11605 = 10'h154 == cnt[9:0] ? $signed(-32'shdd2d) : $signed(_GEN_11604); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11606 = 10'h155 == cnt[9:0] ? $signed(-32'shdd92) : $signed(_GEN_11605); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11607 = 10'h156 == cnt[9:0] ? $signed(-32'shddf7) : $signed(_GEN_11606); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11608 = 10'h157 == cnt[9:0] ? $signed(-32'shde5b) : $signed(_GEN_11607); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11609 = 10'h158 == cnt[9:0] ? $signed(-32'shdebe) : $signed(_GEN_11608); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11610 = 10'h159 == cnt[9:0] ? $signed(-32'shdf21) : $signed(_GEN_11609); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11611 = 10'h15a == cnt[9:0] ? $signed(-32'shdf83) : $signed(_GEN_11610); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11612 = 10'h15b == cnt[9:0] ? $signed(-32'shdfe5) : $signed(_GEN_11611); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11613 = 10'h15c == cnt[9:0] ? $signed(-32'she046) : $signed(_GEN_11612); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11614 = 10'h15d == cnt[9:0] ? $signed(-32'she0a7) : $signed(_GEN_11613); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11615 = 10'h15e == cnt[9:0] ? $signed(-32'she107) : $signed(_GEN_11614); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11616 = 10'h15f == cnt[9:0] ? $signed(-32'she167) : $signed(_GEN_11615); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11617 = 10'h160 == cnt[9:0] ? $signed(-32'she1c6) : $signed(_GEN_11616); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11618 = 10'h161 == cnt[9:0] ? $signed(-32'she224) : $signed(_GEN_11617); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11619 = 10'h162 == cnt[9:0] ? $signed(-32'she282) : $signed(_GEN_11618); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11620 = 10'h163 == cnt[9:0] ? $signed(-32'she2df) : $signed(_GEN_11619); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11621 = 10'h164 == cnt[9:0] ? $signed(-32'she33c) : $signed(_GEN_11620); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11622 = 10'h165 == cnt[9:0] ? $signed(-32'she399) : $signed(_GEN_11621); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11623 = 10'h166 == cnt[9:0] ? $signed(-32'she3f4) : $signed(_GEN_11622); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11624 = 10'h167 == cnt[9:0] ? $signed(-32'she450) : $signed(_GEN_11623); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11625 = 10'h168 == cnt[9:0] ? $signed(-32'she4aa) : $signed(_GEN_11624); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11626 = 10'h169 == cnt[9:0] ? $signed(-32'she504) : $signed(_GEN_11625); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11627 = 10'h16a == cnt[9:0] ? $signed(-32'she55e) : $signed(_GEN_11626); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11628 = 10'h16b == cnt[9:0] ? $signed(-32'she5b7) : $signed(_GEN_11627); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11629 = 10'h16c == cnt[9:0] ? $signed(-32'she610) : $signed(_GEN_11628); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11630 = 10'h16d == cnt[9:0] ? $signed(-32'she667) : $signed(_GEN_11629); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11631 = 10'h16e == cnt[9:0] ? $signed(-32'she6bf) : $signed(_GEN_11630); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11632 = 10'h16f == cnt[9:0] ? $signed(-32'she716) : $signed(_GEN_11631); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11633 = 10'h170 == cnt[9:0] ? $signed(-32'she76c) : $signed(_GEN_11632); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11634 = 10'h171 == cnt[9:0] ? $signed(-32'she7c2) : $signed(_GEN_11633); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11635 = 10'h172 == cnt[9:0] ? $signed(-32'she817) : $signed(_GEN_11634); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11636 = 10'h173 == cnt[9:0] ? $signed(-32'she86b) : $signed(_GEN_11635); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11637 = 10'h174 == cnt[9:0] ? $signed(-32'she8bf) : $signed(_GEN_11636); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11638 = 10'h175 == cnt[9:0] ? $signed(-32'she913) : $signed(_GEN_11637); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11639 = 10'h176 == cnt[9:0] ? $signed(-32'she966) : $signed(_GEN_11638); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11640 = 10'h177 == cnt[9:0] ? $signed(-32'she9b8) : $signed(_GEN_11639); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11641 = 10'h178 == cnt[9:0] ? $signed(-32'shea0a) : $signed(_GEN_11640); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11642 = 10'h179 == cnt[9:0] ? $signed(-32'shea5b) : $signed(_GEN_11641); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11643 = 10'h17a == cnt[9:0] ? $signed(-32'sheaab) : $signed(_GEN_11642); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11644 = 10'h17b == cnt[9:0] ? $signed(-32'sheafc) : $signed(_GEN_11643); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11645 = 10'h17c == cnt[9:0] ? $signed(-32'sheb4b) : $signed(_GEN_11644); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11646 = 10'h17d == cnt[9:0] ? $signed(-32'sheb9a) : $signed(_GEN_11645); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11647 = 10'h17e == cnt[9:0] ? $signed(-32'shebe8) : $signed(_GEN_11646); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11648 = 10'h17f == cnt[9:0] ? $signed(-32'shec36) : $signed(_GEN_11647); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11649 = 10'h180 == cnt[9:0] ? $signed(-32'shec83) : $signed(_GEN_11648); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11650 = 10'h181 == cnt[9:0] ? $signed(-32'shecd0) : $signed(_GEN_11649); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11651 = 10'h182 == cnt[9:0] ? $signed(-32'shed1c) : $signed(_GEN_11650); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11652 = 10'h183 == cnt[9:0] ? $signed(-32'shed68) : $signed(_GEN_11651); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11653 = 10'h184 == cnt[9:0] ? $signed(-32'shedb3) : $signed(_GEN_11652); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11654 = 10'h185 == cnt[9:0] ? $signed(-32'shedfd) : $signed(_GEN_11653); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11655 = 10'h186 == cnt[9:0] ? $signed(-32'shee47) : $signed(_GEN_11654); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11656 = 10'h187 == cnt[9:0] ? $signed(-32'shee90) : $signed(_GEN_11655); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11657 = 10'h188 == cnt[9:0] ? $signed(-32'sheed9) : $signed(_GEN_11656); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11658 = 10'h189 == cnt[9:0] ? $signed(-32'shef21) : $signed(_GEN_11657); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11659 = 10'h18a == cnt[9:0] ? $signed(-32'shef68) : $signed(_GEN_11658); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11660 = 10'h18b == cnt[9:0] ? $signed(-32'shefaf) : $signed(_GEN_11659); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11661 = 10'h18c == cnt[9:0] ? $signed(-32'sheff5) : $signed(_GEN_11660); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11662 = 10'h18d == cnt[9:0] ? $signed(-32'shf03b) : $signed(_GEN_11661); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11663 = 10'h18e == cnt[9:0] ? $signed(-32'shf080) : $signed(_GEN_11662); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11664 = 10'h18f == cnt[9:0] ? $signed(-32'shf0c5) : $signed(_GEN_11663); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11665 = 10'h190 == cnt[9:0] ? $signed(-32'shf109) : $signed(_GEN_11664); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11666 = 10'h191 == cnt[9:0] ? $signed(-32'shf14c) : $signed(_GEN_11665); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11667 = 10'h192 == cnt[9:0] ? $signed(-32'shf18f) : $signed(_GEN_11666); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11668 = 10'h193 == cnt[9:0] ? $signed(-32'shf1d2) : $signed(_GEN_11667); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11669 = 10'h194 == cnt[9:0] ? $signed(-32'shf213) : $signed(_GEN_11668); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11670 = 10'h195 == cnt[9:0] ? $signed(-32'shf254) : $signed(_GEN_11669); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11671 = 10'h196 == cnt[9:0] ? $signed(-32'shf295) : $signed(_GEN_11670); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11672 = 10'h197 == cnt[9:0] ? $signed(-32'shf2d5) : $signed(_GEN_11671); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11673 = 10'h198 == cnt[9:0] ? $signed(-32'shf314) : $signed(_GEN_11672); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11674 = 10'h199 == cnt[9:0] ? $signed(-32'shf353) : $signed(_GEN_11673); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11675 = 10'h19a == cnt[9:0] ? $signed(-32'shf391) : $signed(_GEN_11674); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11676 = 10'h19b == cnt[9:0] ? $signed(-32'shf3cf) : $signed(_GEN_11675); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11677 = 10'h19c == cnt[9:0] ? $signed(-32'shf40c) : $signed(_GEN_11676); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11678 = 10'h19d == cnt[9:0] ? $signed(-32'shf448) : $signed(_GEN_11677); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11679 = 10'h19e == cnt[9:0] ? $signed(-32'shf484) : $signed(_GEN_11678); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11680 = 10'h19f == cnt[9:0] ? $signed(-32'shf4bf) : $signed(_GEN_11679); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11681 = 10'h1a0 == cnt[9:0] ? $signed(-32'shf4fa) : $signed(_GEN_11680); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11682 = 10'h1a1 == cnt[9:0] ? $signed(-32'shf534) : $signed(_GEN_11681); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11683 = 10'h1a2 == cnt[9:0] ? $signed(-32'shf56e) : $signed(_GEN_11682); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11684 = 10'h1a3 == cnt[9:0] ? $signed(-32'shf5a6) : $signed(_GEN_11683); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11685 = 10'h1a4 == cnt[9:0] ? $signed(-32'shf5df) : $signed(_GEN_11684); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11686 = 10'h1a5 == cnt[9:0] ? $signed(-32'shf616) : $signed(_GEN_11685); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11687 = 10'h1a6 == cnt[9:0] ? $signed(-32'shf64e) : $signed(_GEN_11686); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11688 = 10'h1a7 == cnt[9:0] ? $signed(-32'shf684) : $signed(_GEN_11687); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11689 = 10'h1a8 == cnt[9:0] ? $signed(-32'shf6ba) : $signed(_GEN_11688); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11690 = 10'h1a9 == cnt[9:0] ? $signed(-32'shf6ef) : $signed(_GEN_11689); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11691 = 10'h1aa == cnt[9:0] ? $signed(-32'shf724) : $signed(_GEN_11690); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11692 = 10'h1ab == cnt[9:0] ? $signed(-32'shf758) : $signed(_GEN_11691); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11693 = 10'h1ac == cnt[9:0] ? $signed(-32'shf78c) : $signed(_GEN_11692); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11694 = 10'h1ad == cnt[9:0] ? $signed(-32'shf7bf) : $signed(_GEN_11693); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11695 = 10'h1ae == cnt[9:0] ? $signed(-32'shf7f1) : $signed(_GEN_11694); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11696 = 10'h1af == cnt[9:0] ? $signed(-32'shf823) : $signed(_GEN_11695); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11697 = 10'h1b0 == cnt[9:0] ? $signed(-32'shf854) : $signed(_GEN_11696); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11698 = 10'h1b1 == cnt[9:0] ? $signed(-32'shf885) : $signed(_GEN_11697); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11699 = 10'h1b2 == cnt[9:0] ? $signed(-32'shf8b4) : $signed(_GEN_11698); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11700 = 10'h1b3 == cnt[9:0] ? $signed(-32'shf8e4) : $signed(_GEN_11699); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11701 = 10'h1b4 == cnt[9:0] ? $signed(-32'shf913) : $signed(_GEN_11700); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11702 = 10'h1b5 == cnt[9:0] ? $signed(-32'shf941) : $signed(_GEN_11701); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11703 = 10'h1b6 == cnt[9:0] ? $signed(-32'shf96e) : $signed(_GEN_11702); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11704 = 10'h1b7 == cnt[9:0] ? $signed(-32'shf99b) : $signed(_GEN_11703); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11705 = 10'h1b8 == cnt[9:0] ? $signed(-32'shf9c8) : $signed(_GEN_11704); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11706 = 10'h1b9 == cnt[9:0] ? $signed(-32'shf9f3) : $signed(_GEN_11705); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11707 = 10'h1ba == cnt[9:0] ? $signed(-32'shfa1f) : $signed(_GEN_11706); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11708 = 10'h1bb == cnt[9:0] ? $signed(-32'shfa49) : $signed(_GEN_11707); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11709 = 10'h1bc == cnt[9:0] ? $signed(-32'shfa73) : $signed(_GEN_11708); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11710 = 10'h1bd == cnt[9:0] ? $signed(-32'shfa9c) : $signed(_GEN_11709); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11711 = 10'h1be == cnt[9:0] ? $signed(-32'shfac5) : $signed(_GEN_11710); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11712 = 10'h1bf == cnt[9:0] ? $signed(-32'shfaed) : $signed(_GEN_11711); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11713 = 10'h1c0 == cnt[9:0] ? $signed(-32'shfb15) : $signed(_GEN_11712); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11714 = 10'h1c1 == cnt[9:0] ? $signed(-32'shfb3c) : $signed(_GEN_11713); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11715 = 10'h1c2 == cnt[9:0] ? $signed(-32'shfb62) : $signed(_GEN_11714); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11716 = 10'h1c3 == cnt[9:0] ? $signed(-32'shfb88) : $signed(_GEN_11715); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11717 = 10'h1c4 == cnt[9:0] ? $signed(-32'shfbad) : $signed(_GEN_11716); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11718 = 10'h1c5 == cnt[9:0] ? $signed(-32'shfbd1) : $signed(_GEN_11717); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11719 = 10'h1c6 == cnt[9:0] ? $signed(-32'shfbf5) : $signed(_GEN_11718); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11720 = 10'h1c7 == cnt[9:0] ? $signed(-32'shfc18) : $signed(_GEN_11719); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11721 = 10'h1c8 == cnt[9:0] ? $signed(-32'shfc3b) : $signed(_GEN_11720); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11722 = 10'h1c9 == cnt[9:0] ? $signed(-32'shfc5d) : $signed(_GEN_11721); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11723 = 10'h1ca == cnt[9:0] ? $signed(-32'shfc7f) : $signed(_GEN_11722); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11724 = 10'h1cb == cnt[9:0] ? $signed(-32'shfca0) : $signed(_GEN_11723); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11725 = 10'h1cc == cnt[9:0] ? $signed(-32'shfcc0) : $signed(_GEN_11724); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11726 = 10'h1cd == cnt[9:0] ? $signed(-32'shfcdf) : $signed(_GEN_11725); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11727 = 10'h1ce == cnt[9:0] ? $signed(-32'shfcfe) : $signed(_GEN_11726); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11728 = 10'h1cf == cnt[9:0] ? $signed(-32'shfd1d) : $signed(_GEN_11727); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11729 = 10'h1d0 == cnt[9:0] ? $signed(-32'shfd3b) : $signed(_GEN_11728); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11730 = 10'h1d1 == cnt[9:0] ? $signed(-32'shfd58) : $signed(_GEN_11729); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11731 = 10'h1d2 == cnt[9:0] ? $signed(-32'shfd74) : $signed(_GEN_11730); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11732 = 10'h1d3 == cnt[9:0] ? $signed(-32'shfd90) : $signed(_GEN_11731); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11733 = 10'h1d4 == cnt[9:0] ? $signed(-32'shfdac) : $signed(_GEN_11732); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11734 = 10'h1d5 == cnt[9:0] ? $signed(-32'shfdc7) : $signed(_GEN_11733); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11735 = 10'h1d6 == cnt[9:0] ? $signed(-32'shfde1) : $signed(_GEN_11734); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11736 = 10'h1d7 == cnt[9:0] ? $signed(-32'shfdfa) : $signed(_GEN_11735); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11737 = 10'h1d8 == cnt[9:0] ? $signed(-32'shfe13) : $signed(_GEN_11736); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11738 = 10'h1d9 == cnt[9:0] ? $signed(-32'shfe2b) : $signed(_GEN_11737); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11739 = 10'h1da == cnt[9:0] ? $signed(-32'shfe43) : $signed(_GEN_11738); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11740 = 10'h1db == cnt[9:0] ? $signed(-32'shfe5a) : $signed(_GEN_11739); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11741 = 10'h1dc == cnt[9:0] ? $signed(-32'shfe71) : $signed(_GEN_11740); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11742 = 10'h1dd == cnt[9:0] ? $signed(-32'shfe87) : $signed(_GEN_11741); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11743 = 10'h1de == cnt[9:0] ? $signed(-32'shfe9c) : $signed(_GEN_11742); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11744 = 10'h1df == cnt[9:0] ? $signed(-32'shfeb0) : $signed(_GEN_11743); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11745 = 10'h1e0 == cnt[9:0] ? $signed(-32'shfec4) : $signed(_GEN_11744); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11746 = 10'h1e1 == cnt[9:0] ? $signed(-32'shfed8) : $signed(_GEN_11745); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11747 = 10'h1e2 == cnt[9:0] ? $signed(-32'shfeeb) : $signed(_GEN_11746); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11748 = 10'h1e3 == cnt[9:0] ? $signed(-32'shfefd) : $signed(_GEN_11747); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11749 = 10'h1e4 == cnt[9:0] ? $signed(-32'shff0e) : $signed(_GEN_11748); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11750 = 10'h1e5 == cnt[9:0] ? $signed(-32'shff1f) : $signed(_GEN_11749); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11751 = 10'h1e6 == cnt[9:0] ? $signed(-32'shff30) : $signed(_GEN_11750); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11752 = 10'h1e7 == cnt[9:0] ? $signed(-32'shff3f) : $signed(_GEN_11751); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11753 = 10'h1e8 == cnt[9:0] ? $signed(-32'shff4e) : $signed(_GEN_11752); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11754 = 10'h1e9 == cnt[9:0] ? $signed(-32'shff5d) : $signed(_GEN_11753); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11755 = 10'h1ea == cnt[9:0] ? $signed(-32'shff6b) : $signed(_GEN_11754); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11756 = 10'h1eb == cnt[9:0] ? $signed(-32'shff78) : $signed(_GEN_11755); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11757 = 10'h1ec == cnt[9:0] ? $signed(-32'shff85) : $signed(_GEN_11756); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11758 = 10'h1ed == cnt[9:0] ? $signed(-32'shff91) : $signed(_GEN_11757); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11759 = 10'h1ee == cnt[9:0] ? $signed(-32'shff9c) : $signed(_GEN_11758); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11760 = 10'h1ef == cnt[9:0] ? $signed(-32'shffa7) : $signed(_GEN_11759); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11761 = 10'h1f0 == cnt[9:0] ? $signed(-32'shffb1) : $signed(_GEN_11760); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11762 = 10'h1f1 == cnt[9:0] ? $signed(-32'shffbb) : $signed(_GEN_11761); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11763 = 10'h1f2 == cnt[9:0] ? $signed(-32'shffc4) : $signed(_GEN_11762); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11764 = 10'h1f3 == cnt[9:0] ? $signed(-32'shffcc) : $signed(_GEN_11763); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11765 = 10'h1f4 == cnt[9:0] ? $signed(-32'shffd4) : $signed(_GEN_11764); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11766 = 10'h1f5 == cnt[9:0] ? $signed(-32'shffdb) : $signed(_GEN_11765); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11767 = 10'h1f6 == cnt[9:0] ? $signed(-32'shffe1) : $signed(_GEN_11766); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11768 = 10'h1f7 == cnt[9:0] ? $signed(-32'shffe7) : $signed(_GEN_11767); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11769 = 10'h1f8 == cnt[9:0] ? $signed(-32'shffec) : $signed(_GEN_11768); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11770 = 10'h1f9 == cnt[9:0] ? $signed(-32'shfff1) : $signed(_GEN_11769); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11771 = 10'h1fa == cnt[9:0] ? $signed(-32'shfff5) : $signed(_GEN_11770); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11772 = 10'h1fb == cnt[9:0] ? $signed(-32'shfff8) : $signed(_GEN_11771); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11773 = 10'h1fc == cnt[9:0] ? $signed(-32'shfffb) : $signed(_GEN_11772); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11774 = 10'h1fd == cnt[9:0] ? $signed(-32'shfffd) : $signed(_GEN_11773); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11775 = 10'h1fe == cnt[9:0] ? $signed(-32'shffff) : $signed(_GEN_11774); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11776 = 10'h1ff == cnt[9:0] ? $signed(-32'sh10000) : $signed(_GEN_11775); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11777 = 10'h200 == cnt[9:0] ? $signed(-32'sh10000) : $signed(_GEN_11776); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11778 = 10'h201 == cnt[9:0] ? $signed(-32'sh10000) : $signed(_GEN_11777); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11779 = 10'h202 == cnt[9:0] ? $signed(-32'shffff) : $signed(_GEN_11778); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11780 = 10'h203 == cnt[9:0] ? $signed(-32'shfffd) : $signed(_GEN_11779); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11781 = 10'h204 == cnt[9:0] ? $signed(-32'shfffb) : $signed(_GEN_11780); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11782 = 10'h205 == cnt[9:0] ? $signed(-32'shfff8) : $signed(_GEN_11781); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11783 = 10'h206 == cnt[9:0] ? $signed(-32'shfff5) : $signed(_GEN_11782); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11784 = 10'h207 == cnt[9:0] ? $signed(-32'shfff1) : $signed(_GEN_11783); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11785 = 10'h208 == cnt[9:0] ? $signed(-32'shffec) : $signed(_GEN_11784); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11786 = 10'h209 == cnt[9:0] ? $signed(-32'shffe7) : $signed(_GEN_11785); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11787 = 10'h20a == cnt[9:0] ? $signed(-32'shffe1) : $signed(_GEN_11786); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11788 = 10'h20b == cnt[9:0] ? $signed(-32'shffdb) : $signed(_GEN_11787); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11789 = 10'h20c == cnt[9:0] ? $signed(-32'shffd4) : $signed(_GEN_11788); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11790 = 10'h20d == cnt[9:0] ? $signed(-32'shffcc) : $signed(_GEN_11789); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11791 = 10'h20e == cnt[9:0] ? $signed(-32'shffc4) : $signed(_GEN_11790); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11792 = 10'h20f == cnt[9:0] ? $signed(-32'shffbb) : $signed(_GEN_11791); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11793 = 10'h210 == cnt[9:0] ? $signed(-32'shffb1) : $signed(_GEN_11792); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11794 = 10'h211 == cnt[9:0] ? $signed(-32'shffa7) : $signed(_GEN_11793); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11795 = 10'h212 == cnt[9:0] ? $signed(-32'shff9c) : $signed(_GEN_11794); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11796 = 10'h213 == cnt[9:0] ? $signed(-32'shff91) : $signed(_GEN_11795); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11797 = 10'h214 == cnt[9:0] ? $signed(-32'shff85) : $signed(_GEN_11796); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11798 = 10'h215 == cnt[9:0] ? $signed(-32'shff78) : $signed(_GEN_11797); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11799 = 10'h216 == cnt[9:0] ? $signed(-32'shff6b) : $signed(_GEN_11798); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11800 = 10'h217 == cnt[9:0] ? $signed(-32'shff5d) : $signed(_GEN_11799); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11801 = 10'h218 == cnt[9:0] ? $signed(-32'shff4e) : $signed(_GEN_11800); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11802 = 10'h219 == cnt[9:0] ? $signed(-32'shff3f) : $signed(_GEN_11801); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11803 = 10'h21a == cnt[9:0] ? $signed(-32'shff30) : $signed(_GEN_11802); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11804 = 10'h21b == cnt[9:0] ? $signed(-32'shff1f) : $signed(_GEN_11803); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11805 = 10'h21c == cnt[9:0] ? $signed(-32'shff0e) : $signed(_GEN_11804); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11806 = 10'h21d == cnt[9:0] ? $signed(-32'shfefd) : $signed(_GEN_11805); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11807 = 10'h21e == cnt[9:0] ? $signed(-32'shfeeb) : $signed(_GEN_11806); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11808 = 10'h21f == cnt[9:0] ? $signed(-32'shfed8) : $signed(_GEN_11807); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11809 = 10'h220 == cnt[9:0] ? $signed(-32'shfec4) : $signed(_GEN_11808); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11810 = 10'h221 == cnt[9:0] ? $signed(-32'shfeb0) : $signed(_GEN_11809); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11811 = 10'h222 == cnt[9:0] ? $signed(-32'shfe9c) : $signed(_GEN_11810); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11812 = 10'h223 == cnt[9:0] ? $signed(-32'shfe87) : $signed(_GEN_11811); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11813 = 10'h224 == cnt[9:0] ? $signed(-32'shfe71) : $signed(_GEN_11812); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11814 = 10'h225 == cnt[9:0] ? $signed(-32'shfe5a) : $signed(_GEN_11813); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11815 = 10'h226 == cnt[9:0] ? $signed(-32'shfe43) : $signed(_GEN_11814); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11816 = 10'h227 == cnt[9:0] ? $signed(-32'shfe2b) : $signed(_GEN_11815); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11817 = 10'h228 == cnt[9:0] ? $signed(-32'shfe13) : $signed(_GEN_11816); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11818 = 10'h229 == cnt[9:0] ? $signed(-32'shfdfa) : $signed(_GEN_11817); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11819 = 10'h22a == cnt[9:0] ? $signed(-32'shfde1) : $signed(_GEN_11818); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11820 = 10'h22b == cnt[9:0] ? $signed(-32'shfdc7) : $signed(_GEN_11819); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11821 = 10'h22c == cnt[9:0] ? $signed(-32'shfdac) : $signed(_GEN_11820); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11822 = 10'h22d == cnt[9:0] ? $signed(-32'shfd90) : $signed(_GEN_11821); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11823 = 10'h22e == cnt[9:0] ? $signed(-32'shfd74) : $signed(_GEN_11822); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11824 = 10'h22f == cnt[9:0] ? $signed(-32'shfd58) : $signed(_GEN_11823); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11825 = 10'h230 == cnt[9:0] ? $signed(-32'shfd3b) : $signed(_GEN_11824); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11826 = 10'h231 == cnt[9:0] ? $signed(-32'shfd1d) : $signed(_GEN_11825); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11827 = 10'h232 == cnt[9:0] ? $signed(-32'shfcfe) : $signed(_GEN_11826); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11828 = 10'h233 == cnt[9:0] ? $signed(-32'shfcdf) : $signed(_GEN_11827); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11829 = 10'h234 == cnt[9:0] ? $signed(-32'shfcc0) : $signed(_GEN_11828); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11830 = 10'h235 == cnt[9:0] ? $signed(-32'shfca0) : $signed(_GEN_11829); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11831 = 10'h236 == cnt[9:0] ? $signed(-32'shfc7f) : $signed(_GEN_11830); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11832 = 10'h237 == cnt[9:0] ? $signed(-32'shfc5d) : $signed(_GEN_11831); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11833 = 10'h238 == cnt[9:0] ? $signed(-32'shfc3b) : $signed(_GEN_11832); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11834 = 10'h239 == cnt[9:0] ? $signed(-32'shfc18) : $signed(_GEN_11833); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11835 = 10'h23a == cnt[9:0] ? $signed(-32'shfbf5) : $signed(_GEN_11834); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11836 = 10'h23b == cnt[9:0] ? $signed(-32'shfbd1) : $signed(_GEN_11835); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11837 = 10'h23c == cnt[9:0] ? $signed(-32'shfbad) : $signed(_GEN_11836); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11838 = 10'h23d == cnt[9:0] ? $signed(-32'shfb88) : $signed(_GEN_11837); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11839 = 10'h23e == cnt[9:0] ? $signed(-32'shfb62) : $signed(_GEN_11838); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11840 = 10'h23f == cnt[9:0] ? $signed(-32'shfb3c) : $signed(_GEN_11839); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11841 = 10'h240 == cnt[9:0] ? $signed(-32'shfb15) : $signed(_GEN_11840); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11842 = 10'h241 == cnt[9:0] ? $signed(-32'shfaed) : $signed(_GEN_11841); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11843 = 10'h242 == cnt[9:0] ? $signed(-32'shfac5) : $signed(_GEN_11842); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11844 = 10'h243 == cnt[9:0] ? $signed(-32'shfa9c) : $signed(_GEN_11843); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11845 = 10'h244 == cnt[9:0] ? $signed(-32'shfa73) : $signed(_GEN_11844); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11846 = 10'h245 == cnt[9:0] ? $signed(-32'shfa49) : $signed(_GEN_11845); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11847 = 10'h246 == cnt[9:0] ? $signed(-32'shfa1f) : $signed(_GEN_11846); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11848 = 10'h247 == cnt[9:0] ? $signed(-32'shf9f3) : $signed(_GEN_11847); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11849 = 10'h248 == cnt[9:0] ? $signed(-32'shf9c8) : $signed(_GEN_11848); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11850 = 10'h249 == cnt[9:0] ? $signed(-32'shf99b) : $signed(_GEN_11849); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11851 = 10'h24a == cnt[9:0] ? $signed(-32'shf96e) : $signed(_GEN_11850); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11852 = 10'h24b == cnt[9:0] ? $signed(-32'shf941) : $signed(_GEN_11851); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11853 = 10'h24c == cnt[9:0] ? $signed(-32'shf913) : $signed(_GEN_11852); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11854 = 10'h24d == cnt[9:0] ? $signed(-32'shf8e4) : $signed(_GEN_11853); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11855 = 10'h24e == cnt[9:0] ? $signed(-32'shf8b4) : $signed(_GEN_11854); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11856 = 10'h24f == cnt[9:0] ? $signed(-32'shf885) : $signed(_GEN_11855); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11857 = 10'h250 == cnt[9:0] ? $signed(-32'shf854) : $signed(_GEN_11856); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11858 = 10'h251 == cnt[9:0] ? $signed(-32'shf823) : $signed(_GEN_11857); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11859 = 10'h252 == cnt[9:0] ? $signed(-32'shf7f1) : $signed(_GEN_11858); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11860 = 10'h253 == cnt[9:0] ? $signed(-32'shf7bf) : $signed(_GEN_11859); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11861 = 10'h254 == cnt[9:0] ? $signed(-32'shf78c) : $signed(_GEN_11860); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11862 = 10'h255 == cnt[9:0] ? $signed(-32'shf758) : $signed(_GEN_11861); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11863 = 10'h256 == cnt[9:0] ? $signed(-32'shf724) : $signed(_GEN_11862); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11864 = 10'h257 == cnt[9:0] ? $signed(-32'shf6ef) : $signed(_GEN_11863); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11865 = 10'h258 == cnt[9:0] ? $signed(-32'shf6ba) : $signed(_GEN_11864); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11866 = 10'h259 == cnt[9:0] ? $signed(-32'shf684) : $signed(_GEN_11865); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11867 = 10'h25a == cnt[9:0] ? $signed(-32'shf64e) : $signed(_GEN_11866); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11868 = 10'h25b == cnt[9:0] ? $signed(-32'shf616) : $signed(_GEN_11867); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11869 = 10'h25c == cnt[9:0] ? $signed(-32'shf5df) : $signed(_GEN_11868); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11870 = 10'h25d == cnt[9:0] ? $signed(-32'shf5a6) : $signed(_GEN_11869); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11871 = 10'h25e == cnt[9:0] ? $signed(-32'shf56e) : $signed(_GEN_11870); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11872 = 10'h25f == cnt[9:0] ? $signed(-32'shf534) : $signed(_GEN_11871); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11873 = 10'h260 == cnt[9:0] ? $signed(-32'shf4fa) : $signed(_GEN_11872); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11874 = 10'h261 == cnt[9:0] ? $signed(-32'shf4bf) : $signed(_GEN_11873); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11875 = 10'h262 == cnt[9:0] ? $signed(-32'shf484) : $signed(_GEN_11874); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11876 = 10'h263 == cnt[9:0] ? $signed(-32'shf448) : $signed(_GEN_11875); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11877 = 10'h264 == cnt[9:0] ? $signed(-32'shf40c) : $signed(_GEN_11876); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11878 = 10'h265 == cnt[9:0] ? $signed(-32'shf3cf) : $signed(_GEN_11877); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11879 = 10'h266 == cnt[9:0] ? $signed(-32'shf391) : $signed(_GEN_11878); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11880 = 10'h267 == cnt[9:0] ? $signed(-32'shf353) : $signed(_GEN_11879); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11881 = 10'h268 == cnt[9:0] ? $signed(-32'shf314) : $signed(_GEN_11880); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11882 = 10'h269 == cnt[9:0] ? $signed(-32'shf2d5) : $signed(_GEN_11881); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11883 = 10'h26a == cnt[9:0] ? $signed(-32'shf295) : $signed(_GEN_11882); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11884 = 10'h26b == cnt[9:0] ? $signed(-32'shf254) : $signed(_GEN_11883); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11885 = 10'h26c == cnt[9:0] ? $signed(-32'shf213) : $signed(_GEN_11884); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11886 = 10'h26d == cnt[9:0] ? $signed(-32'shf1d2) : $signed(_GEN_11885); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11887 = 10'h26e == cnt[9:0] ? $signed(-32'shf18f) : $signed(_GEN_11886); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11888 = 10'h26f == cnt[9:0] ? $signed(-32'shf14c) : $signed(_GEN_11887); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11889 = 10'h270 == cnt[9:0] ? $signed(-32'shf109) : $signed(_GEN_11888); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11890 = 10'h271 == cnt[9:0] ? $signed(-32'shf0c5) : $signed(_GEN_11889); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11891 = 10'h272 == cnt[9:0] ? $signed(-32'shf080) : $signed(_GEN_11890); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11892 = 10'h273 == cnt[9:0] ? $signed(-32'shf03b) : $signed(_GEN_11891); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11893 = 10'h274 == cnt[9:0] ? $signed(-32'sheff5) : $signed(_GEN_11892); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11894 = 10'h275 == cnt[9:0] ? $signed(-32'shefaf) : $signed(_GEN_11893); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11895 = 10'h276 == cnt[9:0] ? $signed(-32'shef68) : $signed(_GEN_11894); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11896 = 10'h277 == cnt[9:0] ? $signed(-32'shef21) : $signed(_GEN_11895); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11897 = 10'h278 == cnt[9:0] ? $signed(-32'sheed9) : $signed(_GEN_11896); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11898 = 10'h279 == cnt[9:0] ? $signed(-32'shee90) : $signed(_GEN_11897); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11899 = 10'h27a == cnt[9:0] ? $signed(-32'shee47) : $signed(_GEN_11898); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11900 = 10'h27b == cnt[9:0] ? $signed(-32'shedfd) : $signed(_GEN_11899); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11901 = 10'h27c == cnt[9:0] ? $signed(-32'shedb3) : $signed(_GEN_11900); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11902 = 10'h27d == cnt[9:0] ? $signed(-32'shed68) : $signed(_GEN_11901); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11903 = 10'h27e == cnt[9:0] ? $signed(-32'shed1c) : $signed(_GEN_11902); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11904 = 10'h27f == cnt[9:0] ? $signed(-32'shecd0) : $signed(_GEN_11903); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11905 = 10'h280 == cnt[9:0] ? $signed(-32'shec83) : $signed(_GEN_11904); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11906 = 10'h281 == cnt[9:0] ? $signed(-32'shec36) : $signed(_GEN_11905); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11907 = 10'h282 == cnt[9:0] ? $signed(-32'shebe8) : $signed(_GEN_11906); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11908 = 10'h283 == cnt[9:0] ? $signed(-32'sheb9a) : $signed(_GEN_11907); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11909 = 10'h284 == cnt[9:0] ? $signed(-32'sheb4b) : $signed(_GEN_11908); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11910 = 10'h285 == cnt[9:0] ? $signed(-32'sheafc) : $signed(_GEN_11909); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11911 = 10'h286 == cnt[9:0] ? $signed(-32'sheaab) : $signed(_GEN_11910); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11912 = 10'h287 == cnt[9:0] ? $signed(-32'shea5b) : $signed(_GEN_11911); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11913 = 10'h288 == cnt[9:0] ? $signed(-32'shea0a) : $signed(_GEN_11912); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11914 = 10'h289 == cnt[9:0] ? $signed(-32'she9b8) : $signed(_GEN_11913); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11915 = 10'h28a == cnt[9:0] ? $signed(-32'she966) : $signed(_GEN_11914); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11916 = 10'h28b == cnt[9:0] ? $signed(-32'she913) : $signed(_GEN_11915); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11917 = 10'h28c == cnt[9:0] ? $signed(-32'she8bf) : $signed(_GEN_11916); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11918 = 10'h28d == cnt[9:0] ? $signed(-32'she86b) : $signed(_GEN_11917); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11919 = 10'h28e == cnt[9:0] ? $signed(-32'she817) : $signed(_GEN_11918); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11920 = 10'h28f == cnt[9:0] ? $signed(-32'she7c2) : $signed(_GEN_11919); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11921 = 10'h290 == cnt[9:0] ? $signed(-32'she76c) : $signed(_GEN_11920); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11922 = 10'h291 == cnt[9:0] ? $signed(-32'she716) : $signed(_GEN_11921); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11923 = 10'h292 == cnt[9:0] ? $signed(-32'she6bf) : $signed(_GEN_11922); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11924 = 10'h293 == cnt[9:0] ? $signed(-32'she667) : $signed(_GEN_11923); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11925 = 10'h294 == cnt[9:0] ? $signed(-32'she610) : $signed(_GEN_11924); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11926 = 10'h295 == cnt[9:0] ? $signed(-32'she5b7) : $signed(_GEN_11925); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11927 = 10'h296 == cnt[9:0] ? $signed(-32'she55e) : $signed(_GEN_11926); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11928 = 10'h297 == cnt[9:0] ? $signed(-32'she504) : $signed(_GEN_11927); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11929 = 10'h298 == cnt[9:0] ? $signed(-32'she4aa) : $signed(_GEN_11928); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11930 = 10'h299 == cnt[9:0] ? $signed(-32'she450) : $signed(_GEN_11929); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11931 = 10'h29a == cnt[9:0] ? $signed(-32'she3f4) : $signed(_GEN_11930); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11932 = 10'h29b == cnt[9:0] ? $signed(-32'she399) : $signed(_GEN_11931); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11933 = 10'h29c == cnt[9:0] ? $signed(-32'she33c) : $signed(_GEN_11932); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11934 = 10'h29d == cnt[9:0] ? $signed(-32'she2df) : $signed(_GEN_11933); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11935 = 10'h29e == cnt[9:0] ? $signed(-32'she282) : $signed(_GEN_11934); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11936 = 10'h29f == cnt[9:0] ? $signed(-32'she224) : $signed(_GEN_11935); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11937 = 10'h2a0 == cnt[9:0] ? $signed(-32'she1c6) : $signed(_GEN_11936); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11938 = 10'h2a1 == cnt[9:0] ? $signed(-32'she167) : $signed(_GEN_11937); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11939 = 10'h2a2 == cnt[9:0] ? $signed(-32'she107) : $signed(_GEN_11938); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11940 = 10'h2a3 == cnt[9:0] ? $signed(-32'she0a7) : $signed(_GEN_11939); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11941 = 10'h2a4 == cnt[9:0] ? $signed(-32'she046) : $signed(_GEN_11940); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11942 = 10'h2a5 == cnt[9:0] ? $signed(-32'shdfe5) : $signed(_GEN_11941); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11943 = 10'h2a6 == cnt[9:0] ? $signed(-32'shdf83) : $signed(_GEN_11942); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11944 = 10'h2a7 == cnt[9:0] ? $signed(-32'shdf21) : $signed(_GEN_11943); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11945 = 10'h2a8 == cnt[9:0] ? $signed(-32'shdebe) : $signed(_GEN_11944); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11946 = 10'h2a9 == cnt[9:0] ? $signed(-32'shde5b) : $signed(_GEN_11945); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11947 = 10'h2aa == cnt[9:0] ? $signed(-32'shddf7) : $signed(_GEN_11946); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11948 = 10'h2ab == cnt[9:0] ? $signed(-32'shdd92) : $signed(_GEN_11947); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11949 = 10'h2ac == cnt[9:0] ? $signed(-32'shdd2d) : $signed(_GEN_11948); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11950 = 10'h2ad == cnt[9:0] ? $signed(-32'shdcc8) : $signed(_GEN_11949); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11951 = 10'h2ae == cnt[9:0] ? $signed(-32'shdc62) : $signed(_GEN_11950); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11952 = 10'h2af == cnt[9:0] ? $signed(-32'shdbfb) : $signed(_GEN_11951); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11953 = 10'h2b0 == cnt[9:0] ? $signed(-32'shdb94) : $signed(_GEN_11952); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11954 = 10'h2b1 == cnt[9:0] ? $signed(-32'shdb2c) : $signed(_GEN_11953); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11955 = 10'h2b2 == cnt[9:0] ? $signed(-32'shdac4) : $signed(_GEN_11954); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11956 = 10'h2b3 == cnt[9:0] ? $signed(-32'shda5c) : $signed(_GEN_11955); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11957 = 10'h2b4 == cnt[9:0] ? $signed(-32'shd9f2) : $signed(_GEN_11956); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11958 = 10'h2b5 == cnt[9:0] ? $signed(-32'shd989) : $signed(_GEN_11957); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11959 = 10'h2b6 == cnt[9:0] ? $signed(-32'shd91e) : $signed(_GEN_11958); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11960 = 10'h2b7 == cnt[9:0] ? $signed(-32'shd8b4) : $signed(_GEN_11959); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11961 = 10'h2b8 == cnt[9:0] ? $signed(-32'shd848) : $signed(_GEN_11960); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11962 = 10'h2b9 == cnt[9:0] ? $signed(-32'shd7dc) : $signed(_GEN_11961); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11963 = 10'h2ba == cnt[9:0] ? $signed(-32'shd770) : $signed(_GEN_11962); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11964 = 10'h2bb == cnt[9:0] ? $signed(-32'shd703) : $signed(_GEN_11963); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11965 = 10'h2bc == cnt[9:0] ? $signed(-32'shd696) : $signed(_GEN_11964); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11966 = 10'h2bd == cnt[9:0] ? $signed(-32'shd628) : $signed(_GEN_11965); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11967 = 10'h2be == cnt[9:0] ? $signed(-32'shd5ba) : $signed(_GEN_11966); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11968 = 10'h2bf == cnt[9:0] ? $signed(-32'shd54b) : $signed(_GEN_11967); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11969 = 10'h2c0 == cnt[9:0] ? $signed(-32'shd4db) : $signed(_GEN_11968); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11970 = 10'h2c1 == cnt[9:0] ? $signed(-32'shd46b) : $signed(_GEN_11969); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11971 = 10'h2c2 == cnt[9:0] ? $signed(-32'shd3fb) : $signed(_GEN_11970); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11972 = 10'h2c3 == cnt[9:0] ? $signed(-32'shd38a) : $signed(_GEN_11971); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11973 = 10'h2c4 == cnt[9:0] ? $signed(-32'shd318) : $signed(_GEN_11972); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11974 = 10'h2c5 == cnt[9:0] ? $signed(-32'shd2a6) : $signed(_GEN_11973); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11975 = 10'h2c6 == cnt[9:0] ? $signed(-32'shd234) : $signed(_GEN_11974); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11976 = 10'h2c7 == cnt[9:0] ? $signed(-32'shd1c1) : $signed(_GEN_11975); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11977 = 10'h2c8 == cnt[9:0] ? $signed(-32'shd14d) : $signed(_GEN_11976); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11978 = 10'h2c9 == cnt[9:0] ? $signed(-32'shd0d9) : $signed(_GEN_11977); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11979 = 10'h2ca == cnt[9:0] ? $signed(-32'shd065) : $signed(_GEN_11978); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11980 = 10'h2cb == cnt[9:0] ? $signed(-32'shcff0) : $signed(_GEN_11979); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11981 = 10'h2cc == cnt[9:0] ? $signed(-32'shcf7a) : $signed(_GEN_11980); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11982 = 10'h2cd == cnt[9:0] ? $signed(-32'shcf04) : $signed(_GEN_11981); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11983 = 10'h2ce == cnt[9:0] ? $signed(-32'shce8e) : $signed(_GEN_11982); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11984 = 10'h2cf == cnt[9:0] ? $signed(-32'shce17) : $signed(_GEN_11983); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11985 = 10'h2d0 == cnt[9:0] ? $signed(-32'shcd9f) : $signed(_GEN_11984); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11986 = 10'h2d1 == cnt[9:0] ? $signed(-32'shcd27) : $signed(_GEN_11985); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11987 = 10'h2d2 == cnt[9:0] ? $signed(-32'shccae) : $signed(_GEN_11986); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11988 = 10'h2d3 == cnt[9:0] ? $signed(-32'shcc35) : $signed(_GEN_11987); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11989 = 10'h2d4 == cnt[9:0] ? $signed(-32'shcbbc) : $signed(_GEN_11988); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11990 = 10'h2d5 == cnt[9:0] ? $signed(-32'shcb42) : $signed(_GEN_11989); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11991 = 10'h2d6 == cnt[9:0] ? $signed(-32'shcac7) : $signed(_GEN_11990); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11992 = 10'h2d7 == cnt[9:0] ? $signed(-32'shca4d) : $signed(_GEN_11991); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11993 = 10'h2d8 == cnt[9:0] ? $signed(-32'shc9d1) : $signed(_GEN_11992); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11994 = 10'h2d9 == cnt[9:0] ? $signed(-32'shc955) : $signed(_GEN_11993); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11995 = 10'h2da == cnt[9:0] ? $signed(-32'shc8d9) : $signed(_GEN_11994); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11996 = 10'h2db == cnt[9:0] ? $signed(-32'shc85c) : $signed(_GEN_11995); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11997 = 10'h2dc == cnt[9:0] ? $signed(-32'shc7de) : $signed(_GEN_11996); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11998 = 10'h2dd == cnt[9:0] ? $signed(-32'shc761) : $signed(_GEN_11997); // @[FFT.scala 35:12]
  wire [31:0] _GEN_11999 = 10'h2de == cnt[9:0] ? $signed(-32'shc6e2) : $signed(_GEN_11998); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12000 = 10'h2df == cnt[9:0] ? $signed(-32'shc663) : $signed(_GEN_11999); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12001 = 10'h2e0 == cnt[9:0] ? $signed(-32'shc5e4) : $signed(_GEN_12000); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12002 = 10'h2e1 == cnt[9:0] ? $signed(-32'shc564) : $signed(_GEN_12001); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12003 = 10'h2e2 == cnt[9:0] ? $signed(-32'shc4e4) : $signed(_GEN_12002); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12004 = 10'h2e3 == cnt[9:0] ? $signed(-32'shc463) : $signed(_GEN_12003); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12005 = 10'h2e4 == cnt[9:0] ? $signed(-32'shc3e2) : $signed(_GEN_12004); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12006 = 10'h2e5 == cnt[9:0] ? $signed(-32'shc360) : $signed(_GEN_12005); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12007 = 10'h2e6 == cnt[9:0] ? $signed(-32'shc2de) : $signed(_GEN_12006); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12008 = 10'h2e7 == cnt[9:0] ? $signed(-32'shc25c) : $signed(_GEN_12007); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12009 = 10'h2e8 == cnt[9:0] ? $signed(-32'shc1d8) : $signed(_GEN_12008); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12010 = 10'h2e9 == cnt[9:0] ? $signed(-32'shc155) : $signed(_GEN_12009); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12011 = 10'h2ea == cnt[9:0] ? $signed(-32'shc0d1) : $signed(_GEN_12010); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12012 = 10'h2eb == cnt[9:0] ? $signed(-32'shc04c) : $signed(_GEN_12011); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12013 = 10'h2ec == cnt[9:0] ? $signed(-32'shbfc7) : $signed(_GEN_12012); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12014 = 10'h2ed == cnt[9:0] ? $signed(-32'shbf42) : $signed(_GEN_12013); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12015 = 10'h2ee == cnt[9:0] ? $signed(-32'shbebc) : $signed(_GEN_12014); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12016 = 10'h2ef == cnt[9:0] ? $signed(-32'shbe36) : $signed(_GEN_12015); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12017 = 10'h2f0 == cnt[9:0] ? $signed(-32'shbdaf) : $signed(_GEN_12016); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12018 = 10'h2f1 == cnt[9:0] ? $signed(-32'shbd28) : $signed(_GEN_12017); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12019 = 10'h2f2 == cnt[9:0] ? $signed(-32'shbca0) : $signed(_GEN_12018); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12020 = 10'h2f3 == cnt[9:0] ? $signed(-32'shbc18) : $signed(_GEN_12019); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12021 = 10'h2f4 == cnt[9:0] ? $signed(-32'shbb8f) : $signed(_GEN_12020); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12022 = 10'h2f5 == cnt[9:0] ? $signed(-32'shbb06) : $signed(_GEN_12021); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12023 = 10'h2f6 == cnt[9:0] ? $signed(-32'shba7d) : $signed(_GEN_12022); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12024 = 10'h2f7 == cnt[9:0] ? $signed(-32'shb9f3) : $signed(_GEN_12023); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12025 = 10'h2f8 == cnt[9:0] ? $signed(-32'shb968) : $signed(_GEN_12024); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12026 = 10'h2f9 == cnt[9:0] ? $signed(-32'shb8dd) : $signed(_GEN_12025); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12027 = 10'h2fa == cnt[9:0] ? $signed(-32'shb852) : $signed(_GEN_12026); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12028 = 10'h2fb == cnt[9:0] ? $signed(-32'shb7c6) : $signed(_GEN_12027); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12029 = 10'h2fc == cnt[9:0] ? $signed(-32'shb73a) : $signed(_GEN_12028); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12030 = 10'h2fd == cnt[9:0] ? $signed(-32'shb6ad) : $signed(_GEN_12029); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12031 = 10'h2fe == cnt[9:0] ? $signed(-32'shb620) : $signed(_GEN_12030); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12032 = 10'h2ff == cnt[9:0] ? $signed(-32'shb593) : $signed(_GEN_12031); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12033 = 10'h300 == cnt[9:0] ? $signed(-32'shb505) : $signed(_GEN_12032); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12034 = 10'h301 == cnt[9:0] ? $signed(-32'shb477) : $signed(_GEN_12033); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12035 = 10'h302 == cnt[9:0] ? $signed(-32'shb3e8) : $signed(_GEN_12034); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12036 = 10'h303 == cnt[9:0] ? $signed(-32'shb358) : $signed(_GEN_12035); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12037 = 10'h304 == cnt[9:0] ? $signed(-32'shb2c9) : $signed(_GEN_12036); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12038 = 10'h305 == cnt[9:0] ? $signed(-32'shb239) : $signed(_GEN_12037); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12039 = 10'h306 == cnt[9:0] ? $signed(-32'shb1a8) : $signed(_GEN_12038); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12040 = 10'h307 == cnt[9:0] ? $signed(-32'shb117) : $signed(_GEN_12039); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12041 = 10'h308 == cnt[9:0] ? $signed(-32'shb086) : $signed(_GEN_12040); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12042 = 10'h309 == cnt[9:0] ? $signed(-32'shaff4) : $signed(_GEN_12041); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12043 = 10'h30a == cnt[9:0] ? $signed(-32'shaf62) : $signed(_GEN_12042); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12044 = 10'h30b == cnt[9:0] ? $signed(-32'shaecf) : $signed(_GEN_12043); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12045 = 10'h30c == cnt[9:0] ? $signed(-32'shae3c) : $signed(_GEN_12044); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12046 = 10'h30d == cnt[9:0] ? $signed(-32'shada8) : $signed(_GEN_12045); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12047 = 10'h30e == cnt[9:0] ? $signed(-32'shad14) : $signed(_GEN_12046); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12048 = 10'h30f == cnt[9:0] ? $signed(-32'shac80) : $signed(_GEN_12047); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12049 = 10'h310 == cnt[9:0] ? $signed(-32'shabeb) : $signed(_GEN_12048); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12050 = 10'h311 == cnt[9:0] ? $signed(-32'shab56) : $signed(_GEN_12049); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12051 = 10'h312 == cnt[9:0] ? $signed(-32'shaac1) : $signed(_GEN_12050); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12052 = 10'h313 == cnt[9:0] ? $signed(-32'shaa2a) : $signed(_GEN_12051); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12053 = 10'h314 == cnt[9:0] ? $signed(-32'sha994) : $signed(_GEN_12052); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12054 = 10'h315 == cnt[9:0] ? $signed(-32'sha8fd) : $signed(_GEN_12053); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12055 = 10'h316 == cnt[9:0] ? $signed(-32'sha866) : $signed(_GEN_12054); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12056 = 10'h317 == cnt[9:0] ? $signed(-32'sha7ce) : $signed(_GEN_12055); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12057 = 10'h318 == cnt[9:0] ? $signed(-32'sha736) : $signed(_GEN_12056); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12058 = 10'h319 == cnt[9:0] ? $signed(-32'sha69e) : $signed(_GEN_12057); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12059 = 10'h31a == cnt[9:0] ? $signed(-32'sha605) : $signed(_GEN_12058); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12060 = 10'h31b == cnt[9:0] ? $signed(-32'sha56c) : $signed(_GEN_12059); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12061 = 10'h31c == cnt[9:0] ? $signed(-32'sha4d2) : $signed(_GEN_12060); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12062 = 10'h31d == cnt[9:0] ? $signed(-32'sha438) : $signed(_GEN_12061); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12063 = 10'h31e == cnt[9:0] ? $signed(-32'sha39e) : $signed(_GEN_12062); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12064 = 10'h31f == cnt[9:0] ? $signed(-32'sha303) : $signed(_GEN_12063); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12065 = 10'h320 == cnt[9:0] ? $signed(-32'sha268) : $signed(_GEN_12064); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12066 = 10'h321 == cnt[9:0] ? $signed(-32'sha1cc) : $signed(_GEN_12065); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12067 = 10'h322 == cnt[9:0] ? $signed(-32'sha130) : $signed(_GEN_12066); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12068 = 10'h323 == cnt[9:0] ? $signed(-32'sha094) : $signed(_GEN_12067); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12069 = 10'h324 == cnt[9:0] ? $signed(-32'sh9ff7) : $signed(_GEN_12068); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12070 = 10'h325 == cnt[9:0] ? $signed(-32'sh9f5a) : $signed(_GEN_12069); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12071 = 10'h326 == cnt[9:0] ? $signed(-32'sh9ebc) : $signed(_GEN_12070); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12072 = 10'h327 == cnt[9:0] ? $signed(-32'sh9e1e) : $signed(_GEN_12071); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12073 = 10'h328 == cnt[9:0] ? $signed(-32'sh9d80) : $signed(_GEN_12072); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12074 = 10'h329 == cnt[9:0] ? $signed(-32'sh9ce1) : $signed(_GEN_12073); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12075 = 10'h32a == cnt[9:0] ? $signed(-32'sh9c42) : $signed(_GEN_12074); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12076 = 10'h32b == cnt[9:0] ? $signed(-32'sh9ba3) : $signed(_GEN_12075); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12077 = 10'h32c == cnt[9:0] ? $signed(-32'sh9b03) : $signed(_GEN_12076); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12078 = 10'h32d == cnt[9:0] ? $signed(-32'sh9a63) : $signed(_GEN_12077); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12079 = 10'h32e == cnt[9:0] ? $signed(-32'sh99c2) : $signed(_GEN_12078); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12080 = 10'h32f == cnt[9:0] ? $signed(-32'sh9921) : $signed(_GEN_12079); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12081 = 10'h330 == cnt[9:0] ? $signed(-32'sh9880) : $signed(_GEN_12080); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12082 = 10'h331 == cnt[9:0] ? $signed(-32'sh97de) : $signed(_GEN_12081); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12083 = 10'h332 == cnt[9:0] ? $signed(-32'sh973c) : $signed(_GEN_12082); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12084 = 10'h333 == cnt[9:0] ? $signed(-32'sh969a) : $signed(_GEN_12083); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12085 = 10'h334 == cnt[9:0] ? $signed(-32'sh95f7) : $signed(_GEN_12084); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12086 = 10'h335 == cnt[9:0] ? $signed(-32'sh9554) : $signed(_GEN_12085); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12087 = 10'h336 == cnt[9:0] ? $signed(-32'sh94b0) : $signed(_GEN_12086); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12088 = 10'h337 == cnt[9:0] ? $signed(-32'sh940c) : $signed(_GEN_12087); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12089 = 10'h338 == cnt[9:0] ? $signed(-32'sh9368) : $signed(_GEN_12088); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12090 = 10'h339 == cnt[9:0] ? $signed(-32'sh92c4) : $signed(_GEN_12089); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12091 = 10'h33a == cnt[9:0] ? $signed(-32'sh921f) : $signed(_GEN_12090); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12092 = 10'h33b == cnt[9:0] ? $signed(-32'sh9179) : $signed(_GEN_12091); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12093 = 10'h33c == cnt[9:0] ? $signed(-32'sh90d4) : $signed(_GEN_12092); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12094 = 10'h33d == cnt[9:0] ? $signed(-32'sh902e) : $signed(_GEN_12093); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12095 = 10'h33e == cnt[9:0] ? $signed(-32'sh8f88) : $signed(_GEN_12094); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12096 = 10'h33f == cnt[9:0] ? $signed(-32'sh8ee1) : $signed(_GEN_12095); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12097 = 10'h340 == cnt[9:0] ? $signed(-32'sh8e3a) : $signed(_GEN_12096); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12098 = 10'h341 == cnt[9:0] ? $signed(-32'sh8d93) : $signed(_GEN_12097); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12099 = 10'h342 == cnt[9:0] ? $signed(-32'sh8ceb) : $signed(_GEN_12098); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12100 = 10'h343 == cnt[9:0] ? $signed(-32'sh8c43) : $signed(_GEN_12099); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12101 = 10'h344 == cnt[9:0] ? $signed(-32'sh8b9a) : $signed(_GEN_12100); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12102 = 10'h345 == cnt[9:0] ? $signed(-32'sh8af2) : $signed(_GEN_12101); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12103 = 10'h346 == cnt[9:0] ? $signed(-32'sh8a49) : $signed(_GEN_12102); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12104 = 10'h347 == cnt[9:0] ? $signed(-32'sh899f) : $signed(_GEN_12103); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12105 = 10'h348 == cnt[9:0] ? $signed(-32'sh88f6) : $signed(_GEN_12104); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12106 = 10'h349 == cnt[9:0] ? $signed(-32'sh884c) : $signed(_GEN_12105); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12107 = 10'h34a == cnt[9:0] ? $signed(-32'sh87a1) : $signed(_GEN_12106); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12108 = 10'h34b == cnt[9:0] ? $signed(-32'sh86f7) : $signed(_GEN_12107); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12109 = 10'h34c == cnt[9:0] ? $signed(-32'sh864c) : $signed(_GEN_12108); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12110 = 10'h34d == cnt[9:0] ? $signed(-32'sh85a0) : $signed(_GEN_12109); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12111 = 10'h34e == cnt[9:0] ? $signed(-32'sh84f5) : $signed(_GEN_12110); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12112 = 10'h34f == cnt[9:0] ? $signed(-32'sh8449) : $signed(_GEN_12111); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12113 = 10'h350 == cnt[9:0] ? $signed(-32'sh839c) : $signed(_GEN_12112); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12114 = 10'h351 == cnt[9:0] ? $signed(-32'sh82f0) : $signed(_GEN_12113); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12115 = 10'h352 == cnt[9:0] ? $signed(-32'sh8243) : $signed(_GEN_12114); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12116 = 10'h353 == cnt[9:0] ? $signed(-32'sh8195) : $signed(_GEN_12115); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12117 = 10'h354 == cnt[9:0] ? $signed(-32'sh80e8) : $signed(_GEN_12116); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12118 = 10'h355 == cnt[9:0] ? $signed(-32'sh803a) : $signed(_GEN_12117); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12119 = 10'h356 == cnt[9:0] ? $signed(-32'sh7f8c) : $signed(_GEN_12118); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12120 = 10'h357 == cnt[9:0] ? $signed(-32'sh7edd) : $signed(_GEN_12119); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12121 = 10'h358 == cnt[9:0] ? $signed(-32'sh7e2f) : $signed(_GEN_12120); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12122 = 10'h359 == cnt[9:0] ? $signed(-32'sh7d7f) : $signed(_GEN_12121); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12123 = 10'h35a == cnt[9:0] ? $signed(-32'sh7cd0) : $signed(_GEN_12122); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12124 = 10'h35b == cnt[9:0] ? $signed(-32'sh7c20) : $signed(_GEN_12123); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12125 = 10'h35c == cnt[9:0] ? $signed(-32'sh7b70) : $signed(_GEN_12124); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12126 = 10'h35d == cnt[9:0] ? $signed(-32'sh7ac0) : $signed(_GEN_12125); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12127 = 10'h35e == cnt[9:0] ? $signed(-32'sh7a10) : $signed(_GEN_12126); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12128 = 10'h35f == cnt[9:0] ? $signed(-32'sh795f) : $signed(_GEN_12127); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12129 = 10'h360 == cnt[9:0] ? $signed(-32'sh78ad) : $signed(_GEN_12128); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12130 = 10'h361 == cnt[9:0] ? $signed(-32'sh77fc) : $signed(_GEN_12129); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12131 = 10'h362 == cnt[9:0] ? $signed(-32'sh774a) : $signed(_GEN_12130); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12132 = 10'h363 == cnt[9:0] ? $signed(-32'sh7698) : $signed(_GEN_12131); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12133 = 10'h364 == cnt[9:0] ? $signed(-32'sh75e6) : $signed(_GEN_12132); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12134 = 10'h365 == cnt[9:0] ? $signed(-32'sh7533) : $signed(_GEN_12133); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12135 = 10'h366 == cnt[9:0] ? $signed(-32'sh7480) : $signed(_GEN_12134); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12136 = 10'h367 == cnt[9:0] ? $signed(-32'sh73cd) : $signed(_GEN_12135); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12137 = 10'h368 == cnt[9:0] ? $signed(-32'sh731a) : $signed(_GEN_12136); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12138 = 10'h369 == cnt[9:0] ? $signed(-32'sh7266) : $signed(_GEN_12137); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12139 = 10'h36a == cnt[9:0] ? $signed(-32'sh71b2) : $signed(_GEN_12138); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12140 = 10'h36b == cnt[9:0] ? $signed(-32'sh70fe) : $signed(_GEN_12139); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12141 = 10'h36c == cnt[9:0] ? $signed(-32'sh7049) : $signed(_GEN_12140); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12142 = 10'h36d == cnt[9:0] ? $signed(-32'sh6f94) : $signed(_GEN_12141); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12143 = 10'h36e == cnt[9:0] ? $signed(-32'sh6edf) : $signed(_GEN_12142); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12144 = 10'h36f == cnt[9:0] ? $signed(-32'sh6e2a) : $signed(_GEN_12143); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12145 = 10'h370 == cnt[9:0] ? $signed(-32'sh6d74) : $signed(_GEN_12144); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12146 = 10'h371 == cnt[9:0] ? $signed(-32'sh6cbe) : $signed(_GEN_12145); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12147 = 10'h372 == cnt[9:0] ? $signed(-32'sh6c08) : $signed(_GEN_12146); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12148 = 10'h373 == cnt[9:0] ? $signed(-32'sh6b52) : $signed(_GEN_12147); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12149 = 10'h374 == cnt[9:0] ? $signed(-32'sh6a9b) : $signed(_GEN_12148); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12150 = 10'h375 == cnt[9:0] ? $signed(-32'sh69e4) : $signed(_GEN_12149); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12151 = 10'h376 == cnt[9:0] ? $signed(-32'sh692d) : $signed(_GEN_12150); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12152 = 10'h377 == cnt[9:0] ? $signed(-32'sh6876) : $signed(_GEN_12151); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12153 = 10'h378 == cnt[9:0] ? $signed(-32'sh67be) : $signed(_GEN_12152); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12154 = 10'h379 == cnt[9:0] ? $signed(-32'sh6706) : $signed(_GEN_12153); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12155 = 10'h37a == cnt[9:0] ? $signed(-32'sh664e) : $signed(_GEN_12154); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12156 = 10'h37b == cnt[9:0] ? $signed(-32'sh6595) : $signed(_GEN_12155); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12157 = 10'h37c == cnt[9:0] ? $signed(-32'sh64dd) : $signed(_GEN_12156); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12158 = 10'h37d == cnt[9:0] ? $signed(-32'sh6424) : $signed(_GEN_12157); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12159 = 10'h37e == cnt[9:0] ? $signed(-32'sh636b) : $signed(_GEN_12158); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12160 = 10'h37f == cnt[9:0] ? $signed(-32'sh62b1) : $signed(_GEN_12159); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12161 = 10'h380 == cnt[9:0] ? $signed(-32'sh61f8) : $signed(_GEN_12160); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12162 = 10'h381 == cnt[9:0] ? $signed(-32'sh613e) : $signed(_GEN_12161); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12163 = 10'h382 == cnt[9:0] ? $signed(-32'sh6084) : $signed(_GEN_12162); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12164 = 10'h383 == cnt[9:0] ? $signed(-32'sh5fc9) : $signed(_GEN_12163); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12165 = 10'h384 == cnt[9:0] ? $signed(-32'sh5f0f) : $signed(_GEN_12164); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12166 = 10'h385 == cnt[9:0] ? $signed(-32'sh5e54) : $signed(_GEN_12165); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12167 = 10'h386 == cnt[9:0] ? $signed(-32'sh5d99) : $signed(_GEN_12166); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12168 = 10'h387 == cnt[9:0] ? $signed(-32'sh5cde) : $signed(_GEN_12167); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12169 = 10'h388 == cnt[9:0] ? $signed(-32'sh5c22) : $signed(_GEN_12168); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12170 = 10'h389 == cnt[9:0] ? $signed(-32'sh5b66) : $signed(_GEN_12169); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12171 = 10'h38a == cnt[9:0] ? $signed(-32'sh5aaa) : $signed(_GEN_12170); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12172 = 10'h38b == cnt[9:0] ? $signed(-32'sh59ee) : $signed(_GEN_12171); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12173 = 10'h38c == cnt[9:0] ? $signed(-32'sh5932) : $signed(_GEN_12172); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12174 = 10'h38d == cnt[9:0] ? $signed(-32'sh5875) : $signed(_GEN_12173); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12175 = 10'h38e == cnt[9:0] ? $signed(-32'sh57b9) : $signed(_GEN_12174); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12176 = 10'h38f == cnt[9:0] ? $signed(-32'sh56fc) : $signed(_GEN_12175); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12177 = 10'h390 == cnt[9:0] ? $signed(-32'sh563e) : $signed(_GEN_12176); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12178 = 10'h391 == cnt[9:0] ? $signed(-32'sh5581) : $signed(_GEN_12177); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12179 = 10'h392 == cnt[9:0] ? $signed(-32'sh54c3) : $signed(_GEN_12178); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12180 = 10'h393 == cnt[9:0] ? $signed(-32'sh5406) : $signed(_GEN_12179); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12181 = 10'h394 == cnt[9:0] ? $signed(-32'sh5348) : $signed(_GEN_12180); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12182 = 10'h395 == cnt[9:0] ? $signed(-32'sh5289) : $signed(_GEN_12181); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12183 = 10'h396 == cnt[9:0] ? $signed(-32'sh51cb) : $signed(_GEN_12182); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12184 = 10'h397 == cnt[9:0] ? $signed(-32'sh510c) : $signed(_GEN_12183); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12185 = 10'h398 == cnt[9:0] ? $signed(-32'sh504d) : $signed(_GEN_12184); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12186 = 10'h399 == cnt[9:0] ? $signed(-32'sh4f8e) : $signed(_GEN_12185); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12187 = 10'h39a == cnt[9:0] ? $signed(-32'sh4ecf) : $signed(_GEN_12186); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12188 = 10'h39b == cnt[9:0] ? $signed(-32'sh4e10) : $signed(_GEN_12187); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12189 = 10'h39c == cnt[9:0] ? $signed(-32'sh4d50) : $signed(_GEN_12188); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12190 = 10'h39d == cnt[9:0] ? $signed(-32'sh4c90) : $signed(_GEN_12189); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12191 = 10'h39e == cnt[9:0] ? $signed(-32'sh4bd1) : $signed(_GEN_12190); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12192 = 10'h39f == cnt[9:0] ? $signed(-32'sh4b10) : $signed(_GEN_12191); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12193 = 10'h3a0 == cnt[9:0] ? $signed(-32'sh4a50) : $signed(_GEN_12192); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12194 = 10'h3a1 == cnt[9:0] ? $signed(-32'sh4990) : $signed(_GEN_12193); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12195 = 10'h3a2 == cnt[9:0] ? $signed(-32'sh48cf) : $signed(_GEN_12194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12196 = 10'h3a3 == cnt[9:0] ? $signed(-32'sh480e) : $signed(_GEN_12195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12197 = 10'h3a4 == cnt[9:0] ? $signed(-32'sh474d) : $signed(_GEN_12196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12198 = 10'h3a5 == cnt[9:0] ? $signed(-32'sh468c) : $signed(_GEN_12197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12199 = 10'h3a6 == cnt[9:0] ? $signed(-32'sh45cb) : $signed(_GEN_12198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12200 = 10'h3a7 == cnt[9:0] ? $signed(-32'sh4509) : $signed(_GEN_12199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12201 = 10'h3a8 == cnt[9:0] ? $signed(-32'sh4447) : $signed(_GEN_12200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12202 = 10'h3a9 == cnt[9:0] ? $signed(-32'sh4385) : $signed(_GEN_12201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12203 = 10'h3aa == cnt[9:0] ? $signed(-32'sh42c3) : $signed(_GEN_12202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12204 = 10'h3ab == cnt[9:0] ? $signed(-32'sh4201) : $signed(_GEN_12203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12205 = 10'h3ac == cnt[9:0] ? $signed(-32'sh413f) : $signed(_GEN_12204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12206 = 10'h3ad == cnt[9:0] ? $signed(-32'sh407c) : $signed(_GEN_12205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12207 = 10'h3ae == cnt[9:0] ? $signed(-32'sh3fba) : $signed(_GEN_12206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12208 = 10'h3af == cnt[9:0] ? $signed(-32'sh3ef7) : $signed(_GEN_12207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12209 = 10'h3b0 == cnt[9:0] ? $signed(-32'sh3e34) : $signed(_GEN_12208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12210 = 10'h3b1 == cnt[9:0] ? $signed(-32'sh3d71) : $signed(_GEN_12209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12211 = 10'h3b2 == cnt[9:0] ? $signed(-32'sh3cae) : $signed(_GEN_12210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12212 = 10'h3b3 == cnt[9:0] ? $signed(-32'sh3bea) : $signed(_GEN_12211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12213 = 10'h3b4 == cnt[9:0] ? $signed(-32'sh3b27) : $signed(_GEN_12212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12214 = 10'h3b5 == cnt[9:0] ? $signed(-32'sh3a63) : $signed(_GEN_12213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12215 = 10'h3b6 == cnt[9:0] ? $signed(-32'sh399f) : $signed(_GEN_12214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12216 = 10'h3b7 == cnt[9:0] ? $signed(-32'sh38db) : $signed(_GEN_12215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12217 = 10'h3b8 == cnt[9:0] ? $signed(-32'sh3817) : $signed(_GEN_12216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12218 = 10'h3b9 == cnt[9:0] ? $signed(-32'sh3753) : $signed(_GEN_12217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12219 = 10'h3ba == cnt[9:0] ? $signed(-32'sh368e) : $signed(_GEN_12218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12220 = 10'h3bb == cnt[9:0] ? $signed(-32'sh35ca) : $signed(_GEN_12219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12221 = 10'h3bc == cnt[9:0] ? $signed(-32'sh3505) : $signed(_GEN_12220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12222 = 10'h3bd == cnt[9:0] ? $signed(-32'sh3440) : $signed(_GEN_12221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12223 = 10'h3be == cnt[9:0] ? $signed(-32'sh337c) : $signed(_GEN_12222); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12224 = 10'h3bf == cnt[9:0] ? $signed(-32'sh32b7) : $signed(_GEN_12223); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12225 = 10'h3c0 == cnt[9:0] ? $signed(-32'sh31f1) : $signed(_GEN_12224); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12226 = 10'h3c1 == cnt[9:0] ? $signed(-32'sh312c) : $signed(_GEN_12225); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12227 = 10'h3c2 == cnt[9:0] ? $signed(-32'sh3067) : $signed(_GEN_12226); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12228 = 10'h3c3 == cnt[9:0] ? $signed(-32'sh2fa1) : $signed(_GEN_12227); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12229 = 10'h3c4 == cnt[9:0] ? $signed(-32'sh2edc) : $signed(_GEN_12228); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12230 = 10'h3c5 == cnt[9:0] ? $signed(-32'sh2e16) : $signed(_GEN_12229); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12231 = 10'h3c6 == cnt[9:0] ? $signed(-32'sh2d50) : $signed(_GEN_12230); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12232 = 10'h3c7 == cnt[9:0] ? $signed(-32'sh2c8a) : $signed(_GEN_12231); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12233 = 10'h3c8 == cnt[9:0] ? $signed(-32'sh2bc4) : $signed(_GEN_12232); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12234 = 10'h3c9 == cnt[9:0] ? $signed(-32'sh2afe) : $signed(_GEN_12233); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12235 = 10'h3ca == cnt[9:0] ? $signed(-32'sh2a38) : $signed(_GEN_12234); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12236 = 10'h3cb == cnt[9:0] ? $signed(-32'sh2971) : $signed(_GEN_12235); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12237 = 10'h3cc == cnt[9:0] ? $signed(-32'sh28ab) : $signed(_GEN_12236); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12238 = 10'h3cd == cnt[9:0] ? $signed(-32'sh27e4) : $signed(_GEN_12237); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12239 = 10'h3ce == cnt[9:0] ? $signed(-32'sh271e) : $signed(_GEN_12238); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12240 = 10'h3cf == cnt[9:0] ? $signed(-32'sh2657) : $signed(_GEN_12239); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12241 = 10'h3d0 == cnt[9:0] ? $signed(-32'sh2590) : $signed(_GEN_12240); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12242 = 10'h3d1 == cnt[9:0] ? $signed(-32'sh24c9) : $signed(_GEN_12241); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12243 = 10'h3d2 == cnt[9:0] ? $signed(-32'sh2402) : $signed(_GEN_12242); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12244 = 10'h3d3 == cnt[9:0] ? $signed(-32'sh233b) : $signed(_GEN_12243); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12245 = 10'h3d4 == cnt[9:0] ? $signed(-32'sh2274) : $signed(_GEN_12244); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12246 = 10'h3d5 == cnt[9:0] ? $signed(-32'sh21ad) : $signed(_GEN_12245); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12247 = 10'h3d6 == cnt[9:0] ? $signed(-32'sh20e5) : $signed(_GEN_12246); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12248 = 10'h3d7 == cnt[9:0] ? $signed(-32'sh201e) : $signed(_GEN_12247); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12249 = 10'h3d8 == cnt[9:0] ? $signed(-32'sh1f56) : $signed(_GEN_12248); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12250 = 10'h3d9 == cnt[9:0] ? $signed(-32'sh1e8f) : $signed(_GEN_12249); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12251 = 10'h3da == cnt[9:0] ? $signed(-32'sh1dc7) : $signed(_GEN_12250); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12252 = 10'h3db == cnt[9:0] ? $signed(-32'sh1cff) : $signed(_GEN_12251); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12253 = 10'h3dc == cnt[9:0] ? $signed(-32'sh1c38) : $signed(_GEN_12252); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12254 = 10'h3dd == cnt[9:0] ? $signed(-32'sh1b70) : $signed(_GEN_12253); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12255 = 10'h3de == cnt[9:0] ? $signed(-32'sh1aa8) : $signed(_GEN_12254); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12256 = 10'h3df == cnt[9:0] ? $signed(-32'sh19e0) : $signed(_GEN_12255); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12257 = 10'h3e0 == cnt[9:0] ? $signed(-32'sh1918) : $signed(_GEN_12256); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12258 = 10'h3e1 == cnt[9:0] ? $signed(-32'sh1850) : $signed(_GEN_12257); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12259 = 10'h3e2 == cnt[9:0] ? $signed(-32'sh1787) : $signed(_GEN_12258); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12260 = 10'h3e3 == cnt[9:0] ? $signed(-32'sh16bf) : $signed(_GEN_12259); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12261 = 10'h3e4 == cnt[9:0] ? $signed(-32'sh15f7) : $signed(_GEN_12260); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12262 = 10'h3e5 == cnt[9:0] ? $signed(-32'sh152e) : $signed(_GEN_12261); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12263 = 10'h3e6 == cnt[9:0] ? $signed(-32'sh1466) : $signed(_GEN_12262); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12264 = 10'h3e7 == cnt[9:0] ? $signed(-32'sh139e) : $signed(_GEN_12263); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12265 = 10'h3e8 == cnt[9:0] ? $signed(-32'sh12d5) : $signed(_GEN_12264); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12266 = 10'h3e9 == cnt[9:0] ? $signed(-32'sh120d) : $signed(_GEN_12265); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12267 = 10'h3ea == cnt[9:0] ? $signed(-32'sh1144) : $signed(_GEN_12266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12268 = 10'h3eb == cnt[9:0] ? $signed(-32'sh107b) : $signed(_GEN_12267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12269 = 10'h3ec == cnt[9:0] ? $signed(-32'shfb3) : $signed(_GEN_12268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12270 = 10'h3ed == cnt[9:0] ? $signed(-32'sheea) : $signed(_GEN_12269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12271 = 10'h3ee == cnt[9:0] ? $signed(-32'she21) : $signed(_GEN_12270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12272 = 10'h3ef == cnt[9:0] ? $signed(-32'shd59) : $signed(_GEN_12271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12273 = 10'h3f0 == cnt[9:0] ? $signed(-32'shc90) : $signed(_GEN_12272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12274 = 10'h3f1 == cnt[9:0] ? $signed(-32'shbc7) : $signed(_GEN_12273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12275 = 10'h3f2 == cnt[9:0] ? $signed(-32'shafe) : $signed(_GEN_12274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12276 = 10'h3f3 == cnt[9:0] ? $signed(-32'sha35) : $signed(_GEN_12275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12277 = 10'h3f4 == cnt[9:0] ? $signed(-32'sh96c) : $signed(_GEN_12276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12278 = 10'h3f5 == cnt[9:0] ? $signed(-32'sh8a3) : $signed(_GEN_12277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12279 = 10'h3f6 == cnt[9:0] ? $signed(-32'sh7da) : $signed(_GEN_12278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12280 = 10'h3f7 == cnt[9:0] ? $signed(-32'sh711) : $signed(_GEN_12279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12281 = 10'h3f8 == cnt[9:0] ? $signed(-32'sh648) : $signed(_GEN_12280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12282 = 10'h3f9 == cnt[9:0] ? $signed(-32'sh57f) : $signed(_GEN_12281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12283 = 10'h3fa == cnt[9:0] ? $signed(-32'sh4b6) : $signed(_GEN_12282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12284 = 10'h3fb == cnt[9:0] ? $signed(-32'sh3ed) : $signed(_GEN_12283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12285 = 10'h3fc == cnt[9:0] ? $signed(-32'sh324) : $signed(_GEN_12284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12286 = 10'h3fd == cnt[9:0] ? $signed(-32'sh25b) : $signed(_GEN_12285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_12287 = 10'h3fe == cnt[9:0] ? $signed(-32'sh192) : $signed(_GEN_12286); // @[FFT.scala 35:12]
  reg [31:0] _T_3268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6146;
  reg [31:0] _T_3268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6147;
  reg [31:0] _T_3269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6148;
  reg [31:0] _T_3269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6149;
  reg [31:0] _T_3270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6150;
  reg [31:0] _T_3270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6151;
  reg [31:0] _T_3271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6152;
  reg [31:0] _T_3271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6153;
  reg [31:0] _T_3272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6154;
  reg [31:0] _T_3272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6155;
  reg [31:0] _T_3273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6156;
  reg [31:0] _T_3273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6157;
  reg [31:0] _T_3274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6158;
  reg [31:0] _T_3274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6159;
  reg [31:0] _T_3275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6160;
  reg [31:0] _T_3275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6161;
  reg [31:0] _T_3276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6162;
  reg [31:0] _T_3276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6163;
  reg [31:0] _T_3277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6164;
  reg [31:0] _T_3277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6165;
  reg [31:0] _T_3278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6166;
  reg [31:0] _T_3278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6167;
  reg [31:0] _T_3279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6168;
  reg [31:0] _T_3279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6169;
  reg [31:0] _T_3280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6170;
  reg [31:0] _T_3280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6171;
  reg [31:0] _T_3281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6172;
  reg [31:0] _T_3281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6173;
  reg [31:0] _T_3282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6174;
  reg [31:0] _T_3282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6175;
  reg [31:0] _T_3283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6176;
  reg [31:0] _T_3283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6177;
  reg [31:0] _T_3284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6178;
  reg [31:0] _T_3284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6179;
  reg [31:0] _T_3285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6180;
  reg [31:0] _T_3285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6181;
  reg [31:0] _T_3286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6182;
  reg [31:0] _T_3286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6183;
  reg [31:0] _T_3287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6184;
  reg [31:0] _T_3287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6185;
  reg [31:0] _T_3288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6186;
  reg [31:0] _T_3288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6187;
  reg [31:0] _T_3289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6188;
  reg [31:0] _T_3289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6189;
  reg [31:0] _T_3290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6190;
  reg [31:0] _T_3290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6191;
  reg [31:0] _T_3291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6192;
  reg [31:0] _T_3291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6193;
  reg [31:0] _T_3292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6194;
  reg [31:0] _T_3292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6195;
  reg [31:0] _T_3293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6196;
  reg [31:0] _T_3293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6197;
  reg [31:0] _T_3294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6198;
  reg [31:0] _T_3294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6199;
  reg [31:0] _T_3295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6200;
  reg [31:0] _T_3295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6201;
  reg [31:0] _T_3296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6202;
  reg [31:0] _T_3296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6203;
  reg [31:0] _T_3297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6204;
  reg [31:0] _T_3297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6205;
  reg [31:0] _T_3298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6206;
  reg [31:0] _T_3298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6207;
  reg [31:0] _T_3299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6208;
  reg [31:0] _T_3299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6209;
  reg [31:0] _T_3300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6210;
  reg [31:0] _T_3300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6211;
  reg [31:0] _T_3301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6212;
  reg [31:0] _T_3301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6213;
  reg [31:0] _T_3302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6214;
  reg [31:0] _T_3302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6215;
  reg [31:0] _T_3303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6216;
  reg [31:0] _T_3303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6217;
  reg [31:0] _T_3304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6218;
  reg [31:0] _T_3304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6219;
  reg [31:0] _T_3305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6220;
  reg [31:0] _T_3305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6221;
  reg [31:0] _T_3306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6222;
  reg [31:0] _T_3306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6223;
  reg [31:0] _T_3307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6224;
  reg [31:0] _T_3307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6225;
  reg [31:0] _T_3308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6226;
  reg [31:0] _T_3308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6227;
  reg [31:0] _T_3309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6228;
  reg [31:0] _T_3309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6229;
  reg [31:0] _T_3310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6230;
  reg [31:0] _T_3310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6231;
  reg [31:0] _T_3311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6232;
  reg [31:0] _T_3311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6233;
  reg [31:0] _T_3312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6234;
  reg [31:0] _T_3312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6235;
  reg [31:0] _T_3313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6236;
  reg [31:0] _T_3313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6237;
  reg [31:0] _T_3314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6238;
  reg [31:0] _T_3314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6239;
  reg [31:0] _T_3315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6240;
  reg [31:0] _T_3315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6241;
  reg [31:0] _T_3316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6242;
  reg [31:0] _T_3316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6243;
  reg [31:0] _T_3317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6244;
  reg [31:0] _T_3317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6245;
  reg [31:0] _T_3318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6246;
  reg [31:0] _T_3318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6247;
  reg [31:0] _T_3319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6248;
  reg [31:0] _T_3319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6249;
  reg [31:0] _T_3320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6250;
  reg [31:0] _T_3320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6251;
  reg [31:0] _T_3321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6252;
  reg [31:0] _T_3321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6253;
  reg [31:0] _T_3322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6254;
  reg [31:0] _T_3322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6255;
  reg [31:0] _T_3323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6256;
  reg [31:0] _T_3323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6257;
  reg [31:0] _T_3324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6258;
  reg [31:0] _T_3324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6259;
  reg [31:0] _T_3325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6260;
  reg [31:0] _T_3325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6261;
  reg [31:0] _T_3326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6262;
  reg [31:0] _T_3326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6263;
  reg [31:0] _T_3327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6264;
  reg [31:0] _T_3327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6265;
  reg [31:0] _T_3328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6266;
  reg [31:0] _T_3328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6267;
  reg [31:0] _T_3329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6268;
  reg [31:0] _T_3329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6269;
  reg [31:0] _T_3330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6270;
  reg [31:0] _T_3330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6271;
  reg [31:0] _T_3331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6272;
  reg [31:0] _T_3331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6273;
  reg [31:0] _T_3332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6274;
  reg [31:0] _T_3332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6275;
  reg [31:0] _T_3333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6276;
  reg [31:0] _T_3333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6277;
  reg [31:0] _T_3334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6278;
  reg [31:0] _T_3334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6279;
  reg [31:0] _T_3335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6280;
  reg [31:0] _T_3335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6281;
  reg [31:0] _T_3336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6282;
  reg [31:0] _T_3336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6283;
  reg [31:0] _T_3337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6284;
  reg [31:0] _T_3337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6285;
  reg [31:0] _T_3338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6286;
  reg [31:0] _T_3338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6287;
  reg [31:0] _T_3339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6288;
  reg [31:0] _T_3339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6289;
  reg [31:0] _T_3340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6290;
  reg [31:0] _T_3340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6291;
  reg [31:0] _T_3341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6292;
  reg [31:0] _T_3341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6293;
  reg [31:0] _T_3342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6294;
  reg [31:0] _T_3342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6295;
  reg [31:0] _T_3343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6296;
  reg [31:0] _T_3343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6297;
  reg [31:0] _T_3344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6298;
  reg [31:0] _T_3344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6299;
  reg [31:0] _T_3345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6300;
  reg [31:0] _T_3345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6301;
  reg [31:0] _T_3346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6302;
  reg [31:0] _T_3346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6303;
  reg [31:0] _T_3347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6304;
  reg [31:0] _T_3347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6305;
  reg [31:0] _T_3348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6306;
  reg [31:0] _T_3348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6307;
  reg [31:0] _T_3349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6308;
  reg [31:0] _T_3349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6309;
  reg [31:0] _T_3350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6310;
  reg [31:0] _T_3350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6311;
  reg [31:0] _T_3351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6312;
  reg [31:0] _T_3351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6313;
  reg [31:0] _T_3352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6314;
  reg [31:0] _T_3352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6315;
  reg [31:0] _T_3353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6316;
  reg [31:0] _T_3353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6317;
  reg [31:0] _T_3354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6318;
  reg [31:0] _T_3354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6319;
  reg [31:0] _T_3355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6320;
  reg [31:0] _T_3355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6321;
  reg [31:0] _T_3356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6322;
  reg [31:0] _T_3356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6323;
  reg [31:0] _T_3357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6324;
  reg [31:0] _T_3357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6325;
  reg [31:0] _T_3358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6326;
  reg [31:0] _T_3358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6327;
  reg [31:0] _T_3359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6328;
  reg [31:0] _T_3359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6329;
  reg [31:0] _T_3360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6330;
  reg [31:0] _T_3360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6331;
  reg [31:0] _T_3361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6332;
  reg [31:0] _T_3361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6333;
  reg [31:0] _T_3362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6334;
  reg [31:0] _T_3362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6335;
  reg [31:0] _T_3363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6336;
  reg [31:0] _T_3363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6337;
  reg [31:0] _T_3364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6338;
  reg [31:0] _T_3364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6339;
  reg [31:0] _T_3365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6340;
  reg [31:0] _T_3365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6341;
  reg [31:0] _T_3366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6342;
  reg [31:0] _T_3366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6343;
  reg [31:0] _T_3367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6344;
  reg [31:0] _T_3367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6345;
  reg [31:0] _T_3368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6346;
  reg [31:0] _T_3368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6347;
  reg [31:0] _T_3369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6348;
  reg [31:0] _T_3369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6349;
  reg [31:0] _T_3370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6350;
  reg [31:0] _T_3370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6351;
  reg [31:0] _T_3371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6352;
  reg [31:0] _T_3371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6353;
  reg [31:0] _T_3372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6354;
  reg [31:0] _T_3372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6355;
  reg [31:0] _T_3373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6356;
  reg [31:0] _T_3373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6357;
  reg [31:0] _T_3374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6358;
  reg [31:0] _T_3374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6359;
  reg [31:0] _T_3375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6360;
  reg [31:0] _T_3375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6361;
  reg [31:0] _T_3376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6362;
  reg [31:0] _T_3376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6363;
  reg [31:0] _T_3377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6364;
  reg [31:0] _T_3377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6365;
  reg [31:0] _T_3378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6366;
  reg [31:0] _T_3378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6367;
  reg [31:0] _T_3379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6368;
  reg [31:0] _T_3379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6369;
  reg [31:0] _T_3380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6370;
  reg [31:0] _T_3380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6371;
  reg [31:0] _T_3381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6372;
  reg [31:0] _T_3381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6373;
  reg [31:0] _T_3382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6374;
  reg [31:0] _T_3382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6375;
  reg [31:0] _T_3383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6376;
  reg [31:0] _T_3383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6377;
  reg [31:0] _T_3384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6378;
  reg [31:0] _T_3384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6379;
  reg [31:0] _T_3385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6380;
  reg [31:0] _T_3385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6381;
  reg [31:0] _T_3386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6382;
  reg [31:0] _T_3386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6383;
  reg [31:0] _T_3387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6384;
  reg [31:0] _T_3387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6385;
  reg [31:0] _T_3388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6386;
  reg [31:0] _T_3388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6387;
  reg [31:0] _T_3389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6388;
  reg [31:0] _T_3389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6389;
  reg [31:0] _T_3390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6390;
  reg [31:0] _T_3390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6391;
  reg [31:0] _T_3391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6392;
  reg [31:0] _T_3391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6393;
  reg [31:0] _T_3392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6394;
  reg [31:0] _T_3392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6395;
  reg [31:0] _T_3393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6396;
  reg [31:0] _T_3393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6397;
  reg [31:0] _T_3394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6398;
  reg [31:0] _T_3394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6399;
  reg [31:0] _T_3395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6400;
  reg [31:0] _T_3395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6401;
  reg [31:0] _T_3396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6402;
  reg [31:0] _T_3396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6403;
  reg [31:0] _T_3397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6404;
  reg [31:0] _T_3397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6405;
  reg [31:0] _T_3398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6406;
  reg [31:0] _T_3398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6407;
  reg [31:0] _T_3399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6408;
  reg [31:0] _T_3399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6409;
  reg [31:0] _T_3400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6410;
  reg [31:0] _T_3400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6411;
  reg [31:0] _T_3401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6412;
  reg [31:0] _T_3401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6413;
  reg [31:0] _T_3402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6414;
  reg [31:0] _T_3402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6415;
  reg [31:0] _T_3403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6416;
  reg [31:0] _T_3403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6417;
  reg [31:0] _T_3404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6418;
  reg [31:0] _T_3404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6419;
  reg [31:0] _T_3405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6420;
  reg [31:0] _T_3405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6421;
  reg [31:0] _T_3406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6422;
  reg [31:0] _T_3406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6423;
  reg [31:0] _T_3407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6424;
  reg [31:0] _T_3407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6425;
  reg [31:0] _T_3408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6426;
  reg [31:0] _T_3408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6427;
  reg [31:0] _T_3409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6428;
  reg [31:0] _T_3409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6429;
  reg [31:0] _T_3410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6430;
  reg [31:0] _T_3410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6431;
  reg [31:0] _T_3411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6432;
  reg [31:0] _T_3411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6433;
  reg [31:0] _T_3412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6434;
  reg [31:0] _T_3412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6435;
  reg [31:0] _T_3413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6436;
  reg [31:0] _T_3413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6437;
  reg [31:0] _T_3414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6438;
  reg [31:0] _T_3414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6439;
  reg [31:0] _T_3415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6440;
  reg [31:0] _T_3415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6441;
  reg [31:0] _T_3416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6442;
  reg [31:0] _T_3416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6443;
  reg [31:0] _T_3417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6444;
  reg [31:0] _T_3417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6445;
  reg [31:0] _T_3418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6446;
  reg [31:0] _T_3418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6447;
  reg [31:0] _T_3419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6448;
  reg [31:0] _T_3419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6449;
  reg [31:0] _T_3420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6450;
  reg [31:0] _T_3420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6451;
  reg [31:0] _T_3421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6452;
  reg [31:0] _T_3421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6453;
  reg [31:0] _T_3422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6454;
  reg [31:0] _T_3422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6455;
  reg [31:0] _T_3423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6456;
  reg [31:0] _T_3423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6457;
  reg [31:0] _T_3424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6458;
  reg [31:0] _T_3424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6459;
  reg [31:0] _T_3425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6460;
  reg [31:0] _T_3425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6461;
  reg [31:0] _T_3426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6462;
  reg [31:0] _T_3426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6463;
  reg [31:0] _T_3427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6464;
  reg [31:0] _T_3427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6465;
  reg [31:0] _T_3428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6466;
  reg [31:0] _T_3428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6467;
  reg [31:0] _T_3429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6468;
  reg [31:0] _T_3429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6469;
  reg [31:0] _T_3430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6470;
  reg [31:0] _T_3430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6471;
  reg [31:0] _T_3431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6472;
  reg [31:0] _T_3431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6473;
  reg [31:0] _T_3432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6474;
  reg [31:0] _T_3432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6475;
  reg [31:0] _T_3433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6476;
  reg [31:0] _T_3433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6477;
  reg [31:0] _T_3434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6478;
  reg [31:0] _T_3434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6479;
  reg [31:0] _T_3435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6480;
  reg [31:0] _T_3435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6481;
  reg [31:0] _T_3436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6482;
  reg [31:0] _T_3436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6483;
  reg [31:0] _T_3437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6484;
  reg [31:0] _T_3437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6485;
  reg [31:0] _T_3438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6486;
  reg [31:0] _T_3438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6487;
  reg [31:0] _T_3439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6488;
  reg [31:0] _T_3439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6489;
  reg [31:0] _T_3440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6490;
  reg [31:0] _T_3440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6491;
  reg [31:0] _T_3441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6492;
  reg [31:0] _T_3441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6493;
  reg [31:0] _T_3442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6494;
  reg [31:0] _T_3442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6495;
  reg [31:0] _T_3443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6496;
  reg [31:0] _T_3443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6497;
  reg [31:0] _T_3444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6498;
  reg [31:0] _T_3444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6499;
  reg [31:0] _T_3445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6500;
  reg [31:0] _T_3445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6501;
  reg [31:0] _T_3446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6502;
  reg [31:0] _T_3446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6503;
  reg [31:0] _T_3447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6504;
  reg [31:0] _T_3447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6505;
  reg [31:0] _T_3448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6506;
  reg [31:0] _T_3448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6507;
  reg [31:0] _T_3449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6508;
  reg [31:0] _T_3449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6509;
  reg [31:0] _T_3450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6510;
  reg [31:0] _T_3450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6511;
  reg [31:0] _T_3451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6512;
  reg [31:0] _T_3451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6513;
  reg [31:0] _T_3452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6514;
  reg [31:0] _T_3452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6515;
  reg [31:0] _T_3453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6516;
  reg [31:0] _T_3453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6517;
  reg [31:0] _T_3454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6518;
  reg [31:0] _T_3454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6519;
  reg [31:0] _T_3455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6520;
  reg [31:0] _T_3455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6521;
  reg [31:0] _T_3456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6522;
  reg [31:0] _T_3456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6523;
  reg [31:0] _T_3457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6524;
  reg [31:0] _T_3457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6525;
  reg [31:0] _T_3458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6526;
  reg [31:0] _T_3458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6527;
  reg [31:0] _T_3459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6528;
  reg [31:0] _T_3459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6529;
  reg [31:0] _T_3460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6530;
  reg [31:0] _T_3460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6531;
  reg [31:0] _T_3461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6532;
  reg [31:0] _T_3461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6533;
  reg [31:0] _T_3462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6534;
  reg [31:0] _T_3462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6535;
  reg [31:0] _T_3463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6536;
  reg [31:0] _T_3463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6537;
  reg [31:0] _T_3464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6538;
  reg [31:0] _T_3464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6539;
  reg [31:0] _T_3465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6540;
  reg [31:0] _T_3465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6541;
  reg [31:0] _T_3466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6542;
  reg [31:0] _T_3466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6543;
  reg [31:0] _T_3467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6544;
  reg [31:0] _T_3467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6545;
  reg [31:0] _T_3468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6546;
  reg [31:0] _T_3468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6547;
  reg [31:0] _T_3469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6548;
  reg [31:0] _T_3469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6549;
  reg [31:0] _T_3470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6550;
  reg [31:0] _T_3470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6551;
  reg [31:0] _T_3471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6552;
  reg [31:0] _T_3471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6553;
  reg [31:0] _T_3472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6554;
  reg [31:0] _T_3472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6555;
  reg [31:0] _T_3473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6556;
  reg [31:0] _T_3473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6557;
  reg [31:0] _T_3474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6558;
  reg [31:0] _T_3474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6559;
  reg [31:0] _T_3475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6560;
  reg [31:0] _T_3475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6561;
  reg [31:0] _T_3476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6562;
  reg [31:0] _T_3476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6563;
  reg [31:0] _T_3477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6564;
  reg [31:0] _T_3477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6565;
  reg [31:0] _T_3478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6566;
  reg [31:0] _T_3478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6567;
  reg [31:0] _T_3479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6568;
  reg [31:0] _T_3479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6569;
  reg [31:0] _T_3480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6570;
  reg [31:0] _T_3480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6571;
  reg [31:0] _T_3481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6572;
  reg [31:0] _T_3481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6573;
  reg [31:0] _T_3482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6574;
  reg [31:0] _T_3482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6575;
  reg [31:0] _T_3483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6576;
  reg [31:0] _T_3483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6577;
  reg [31:0] _T_3484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6578;
  reg [31:0] _T_3484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6579;
  reg [31:0] _T_3485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6580;
  reg [31:0] _T_3485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6581;
  reg [31:0] _T_3486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6582;
  reg [31:0] _T_3486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6583;
  reg [31:0] _T_3487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6584;
  reg [31:0] _T_3487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6585;
  reg [31:0] _T_3488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6586;
  reg [31:0] _T_3488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6587;
  reg [31:0] _T_3489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6588;
  reg [31:0] _T_3489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6589;
  reg [31:0] _T_3490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6590;
  reg [31:0] _T_3490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6591;
  reg [31:0] _T_3491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6592;
  reg [31:0] _T_3491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6593;
  reg [31:0] _T_3492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6594;
  reg [31:0] _T_3492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6595;
  reg [31:0] _T_3493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6596;
  reg [31:0] _T_3493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6597;
  reg [31:0] _T_3494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6598;
  reg [31:0] _T_3494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6599;
  reg [31:0] _T_3495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6600;
  reg [31:0] _T_3495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6601;
  reg [31:0] _T_3496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6602;
  reg [31:0] _T_3496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6603;
  reg [31:0] _T_3497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6604;
  reg [31:0] _T_3497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6605;
  reg [31:0] _T_3498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6606;
  reg [31:0] _T_3498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6607;
  reg [31:0] _T_3499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6608;
  reg [31:0] _T_3499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6609;
  reg [31:0] _T_3500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6610;
  reg [31:0] _T_3500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6611;
  reg [31:0] _T_3501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6612;
  reg [31:0] _T_3501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6613;
  reg [31:0] _T_3502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6614;
  reg [31:0] _T_3502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6615;
  reg [31:0] _T_3503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6616;
  reg [31:0] _T_3503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6617;
  reg [31:0] _T_3504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6618;
  reg [31:0] _T_3504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6619;
  reg [31:0] _T_3505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6620;
  reg [31:0] _T_3505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6621;
  reg [31:0] _T_3506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6622;
  reg [31:0] _T_3506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6623;
  reg [31:0] _T_3507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6624;
  reg [31:0] _T_3507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6625;
  reg [31:0] _T_3508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6626;
  reg [31:0] _T_3508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6627;
  reg [31:0] _T_3509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6628;
  reg [31:0] _T_3509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6629;
  reg [31:0] _T_3510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6630;
  reg [31:0] _T_3510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6631;
  reg [31:0] _T_3511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6632;
  reg [31:0] _T_3511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6633;
  reg [31:0] _T_3512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6634;
  reg [31:0] _T_3512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6635;
  reg [31:0] _T_3513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6636;
  reg [31:0] _T_3513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6637;
  reg [31:0] _T_3514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6638;
  reg [31:0] _T_3514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6639;
  reg [31:0] _T_3515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6640;
  reg [31:0] _T_3515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6641;
  reg [31:0] _T_3516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6642;
  reg [31:0] _T_3516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6643;
  reg [31:0] _T_3517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6644;
  reg [31:0] _T_3517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6645;
  reg [31:0] _T_3518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6646;
  reg [31:0] _T_3518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6647;
  reg [31:0] _T_3519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6648;
  reg [31:0] _T_3519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6649;
  reg [31:0] _T_3520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6650;
  reg [31:0] _T_3520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6651;
  reg [31:0] _T_3521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6652;
  reg [31:0] _T_3521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6653;
  reg [31:0] _T_3522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6654;
  reg [31:0] _T_3522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6655;
  reg [31:0] _T_3523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6656;
  reg [31:0] _T_3523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6657;
  reg [31:0] _T_3524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6658;
  reg [31:0] _T_3524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6659;
  reg [31:0] _T_3525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6660;
  reg [31:0] _T_3525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6661;
  reg [31:0] _T_3526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6662;
  reg [31:0] _T_3526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6663;
  reg [31:0] _T_3527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6664;
  reg [31:0] _T_3527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6665;
  reg [31:0] _T_3528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6666;
  reg [31:0] _T_3528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6667;
  reg [31:0] _T_3529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6668;
  reg [31:0] _T_3529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6669;
  reg [31:0] _T_3530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6670;
  reg [31:0] _T_3530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6671;
  reg [31:0] _T_3531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6672;
  reg [31:0] _T_3531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6673;
  reg [31:0] _T_3532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6674;
  reg [31:0] _T_3532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6675;
  reg [31:0] _T_3533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6676;
  reg [31:0] _T_3533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6677;
  reg [31:0] _T_3534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6678;
  reg [31:0] _T_3534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6679;
  reg [31:0] _T_3535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6680;
  reg [31:0] _T_3535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6681;
  reg [31:0] _T_3536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6682;
  reg [31:0] _T_3536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6683;
  reg [31:0] _T_3537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6684;
  reg [31:0] _T_3537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6685;
  reg [31:0] _T_3538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6686;
  reg [31:0] _T_3538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6687;
  reg [31:0] _T_3539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6688;
  reg [31:0] _T_3539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6689;
  reg [31:0] _T_3540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6690;
  reg [31:0] _T_3540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6691;
  reg [31:0] _T_3541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6692;
  reg [31:0] _T_3541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6693;
  reg [31:0] _T_3542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6694;
  reg [31:0] _T_3542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6695;
  reg [31:0] _T_3543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6696;
  reg [31:0] _T_3543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6697;
  reg [31:0] _T_3544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6698;
  reg [31:0] _T_3544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6699;
  reg [31:0] _T_3545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6700;
  reg [31:0] _T_3545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6701;
  reg [31:0] _T_3546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6702;
  reg [31:0] _T_3546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6703;
  reg [31:0] _T_3547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6704;
  reg [31:0] _T_3547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6705;
  reg [31:0] _T_3548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6706;
  reg [31:0] _T_3548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6707;
  reg [31:0] _T_3549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6708;
  reg [31:0] _T_3549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6709;
  reg [31:0] _T_3550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6710;
  reg [31:0] _T_3550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6711;
  reg [31:0] _T_3551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6712;
  reg [31:0] _T_3551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6713;
  reg [31:0] _T_3552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6714;
  reg [31:0] _T_3552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6715;
  reg [31:0] _T_3553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6716;
  reg [31:0] _T_3553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6717;
  reg [31:0] _T_3554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6718;
  reg [31:0] _T_3554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6719;
  reg [31:0] _T_3555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6720;
  reg [31:0] _T_3555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6721;
  reg [31:0] _T_3556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6722;
  reg [31:0] _T_3556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6723;
  reg [31:0] _T_3557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6724;
  reg [31:0] _T_3557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6725;
  reg [31:0] _T_3558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6726;
  reg [31:0] _T_3558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6727;
  reg [31:0] _T_3559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6728;
  reg [31:0] _T_3559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6729;
  reg [31:0] _T_3560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6730;
  reg [31:0] _T_3560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6731;
  reg [31:0] _T_3561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6732;
  reg [31:0] _T_3561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6733;
  reg [31:0] _T_3562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6734;
  reg [31:0] _T_3562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6735;
  reg [31:0] _T_3563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6736;
  reg [31:0] _T_3563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6737;
  reg [31:0] _T_3564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6738;
  reg [31:0] _T_3564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6739;
  reg [31:0] _T_3565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6740;
  reg [31:0] _T_3565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6741;
  reg [31:0] _T_3566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6742;
  reg [31:0] _T_3566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6743;
  reg [31:0] _T_3567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6744;
  reg [31:0] _T_3567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6745;
  reg [31:0] _T_3568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6746;
  reg [31:0] _T_3568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6747;
  reg [31:0] _T_3569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6748;
  reg [31:0] _T_3569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6749;
  reg [31:0] _T_3570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6750;
  reg [31:0] _T_3570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6751;
  reg [31:0] _T_3571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6752;
  reg [31:0] _T_3571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6753;
  reg [31:0] _T_3572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6754;
  reg [31:0] _T_3572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6755;
  reg [31:0] _T_3573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6756;
  reg [31:0] _T_3573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6757;
  reg [31:0] _T_3574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6758;
  reg [31:0] _T_3574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6759;
  reg [31:0] _T_3575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6760;
  reg [31:0] _T_3575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6761;
  reg [31:0] _T_3576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6762;
  reg [31:0] _T_3576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6763;
  reg [31:0] _T_3577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6764;
  reg [31:0] _T_3577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6765;
  reg [31:0] _T_3578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6766;
  reg [31:0] _T_3578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6767;
  reg [31:0] _T_3579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6768;
  reg [31:0] _T_3579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6769;
  reg [31:0] _T_3580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6770;
  reg [31:0] _T_3580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6771;
  reg [31:0] _T_3581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6772;
  reg [31:0] _T_3581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6773;
  reg [31:0] _T_3582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6774;
  reg [31:0] _T_3582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6775;
  reg [31:0] _T_3583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6776;
  reg [31:0] _T_3583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6777;
  reg [31:0] _T_3584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6778;
  reg [31:0] _T_3584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6779;
  reg [31:0] _T_3585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6780;
  reg [31:0] _T_3585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6781;
  reg [31:0] _T_3586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6782;
  reg [31:0] _T_3586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6783;
  reg [31:0] _T_3587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6784;
  reg [31:0] _T_3587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6785;
  reg [31:0] _T_3588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6786;
  reg [31:0] _T_3588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6787;
  reg [31:0] _T_3589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6788;
  reg [31:0] _T_3589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6789;
  reg [31:0] _T_3590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6790;
  reg [31:0] _T_3590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6791;
  reg [31:0] _T_3591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6792;
  reg [31:0] _T_3591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6793;
  reg [31:0] _T_3592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6794;
  reg [31:0] _T_3592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6795;
  reg [31:0] _T_3593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6796;
  reg [31:0] _T_3593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6797;
  reg [31:0] _T_3594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6798;
  reg [31:0] _T_3594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6799;
  reg [31:0] _T_3595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6800;
  reg [31:0] _T_3595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6801;
  reg [31:0] _T_3596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6802;
  reg [31:0] _T_3596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6803;
  reg [31:0] _T_3597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6804;
  reg [31:0] _T_3597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6805;
  reg [31:0] _T_3598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6806;
  reg [31:0] _T_3598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6807;
  reg [31:0] _T_3599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6808;
  reg [31:0] _T_3599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6809;
  reg [31:0] _T_3600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6810;
  reg [31:0] _T_3600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6811;
  reg [31:0] _T_3601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6812;
  reg [31:0] _T_3601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6813;
  reg [31:0] _T_3602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6814;
  reg [31:0] _T_3602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6815;
  reg [31:0] _T_3603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6816;
  reg [31:0] _T_3603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6817;
  reg [31:0] _T_3604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6818;
  reg [31:0] _T_3604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6819;
  reg [31:0] _T_3605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6820;
  reg [31:0] _T_3605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6821;
  reg [31:0] _T_3606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6822;
  reg [31:0] _T_3606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6823;
  reg [31:0] _T_3607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6824;
  reg [31:0] _T_3607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6825;
  reg [31:0] _T_3608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6826;
  reg [31:0] _T_3608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6827;
  reg [31:0] _T_3609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6828;
  reg [31:0] _T_3609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6829;
  reg [31:0] _T_3610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6830;
  reg [31:0] _T_3610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6831;
  reg [31:0] _T_3611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6832;
  reg [31:0] _T_3611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6833;
  reg [31:0] _T_3612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6834;
  reg [31:0] _T_3612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6835;
  reg [31:0] _T_3613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6836;
  reg [31:0] _T_3613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6837;
  reg [31:0] _T_3614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6838;
  reg [31:0] _T_3614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6839;
  reg [31:0] _T_3615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6840;
  reg [31:0] _T_3615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6841;
  reg [31:0] _T_3616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6842;
  reg [31:0] _T_3616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6843;
  reg [31:0] _T_3617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6844;
  reg [31:0] _T_3617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6845;
  reg [31:0] _T_3618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6846;
  reg [31:0] _T_3618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6847;
  reg [31:0] _T_3619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6848;
  reg [31:0] _T_3619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6849;
  reg [31:0] _T_3620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6850;
  reg [31:0] _T_3620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6851;
  reg [31:0] _T_3621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6852;
  reg [31:0] _T_3621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6853;
  reg [31:0] _T_3622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6854;
  reg [31:0] _T_3622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6855;
  reg [31:0] _T_3623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6856;
  reg [31:0] _T_3623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6857;
  reg [31:0] _T_3624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6858;
  reg [31:0] _T_3624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6859;
  reg [31:0] _T_3625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6860;
  reg [31:0] _T_3625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6861;
  reg [31:0] _T_3626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6862;
  reg [31:0] _T_3626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6863;
  reg [31:0] _T_3627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6864;
  reg [31:0] _T_3627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6865;
  reg [31:0] _T_3628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6866;
  reg [31:0] _T_3628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6867;
  reg [31:0] _T_3629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6868;
  reg [31:0] _T_3629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6869;
  reg [31:0] _T_3630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6870;
  reg [31:0] _T_3630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6871;
  reg [31:0] _T_3631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6872;
  reg [31:0] _T_3631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6873;
  reg [31:0] _T_3632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6874;
  reg [31:0] _T_3632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6875;
  reg [31:0] _T_3633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6876;
  reg [31:0] _T_3633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6877;
  reg [31:0] _T_3634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6878;
  reg [31:0] _T_3634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6879;
  reg [31:0] _T_3635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6880;
  reg [31:0] _T_3635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6881;
  reg [31:0] _T_3636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6882;
  reg [31:0] _T_3636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6883;
  reg [31:0] _T_3637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6884;
  reg [31:0] _T_3637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6885;
  reg [31:0] _T_3638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6886;
  reg [31:0] _T_3638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6887;
  reg [31:0] _T_3639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6888;
  reg [31:0] _T_3639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6889;
  reg [31:0] _T_3640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6890;
  reg [31:0] _T_3640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6891;
  reg [31:0] _T_3641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6892;
  reg [31:0] _T_3641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6893;
  reg [31:0] _T_3642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6894;
  reg [31:0] _T_3642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6895;
  reg [31:0] _T_3643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6896;
  reg [31:0] _T_3643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6897;
  reg [31:0] _T_3644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6898;
  reg [31:0] _T_3644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6899;
  reg [31:0] _T_3645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6900;
  reg [31:0] _T_3645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6901;
  reg [31:0] _T_3646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6902;
  reg [31:0] _T_3646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6903;
  reg [31:0] _T_3647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6904;
  reg [31:0] _T_3647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6905;
  reg [31:0] _T_3648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6906;
  reg [31:0] _T_3648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6907;
  reg [31:0] _T_3649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6908;
  reg [31:0] _T_3649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6909;
  reg [31:0] _T_3650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6910;
  reg [31:0] _T_3650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6911;
  reg [31:0] _T_3651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6912;
  reg [31:0] _T_3651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6913;
  reg [31:0] _T_3652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6914;
  reg [31:0] _T_3652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6915;
  reg [31:0] _T_3653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6916;
  reg [31:0] _T_3653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6917;
  reg [31:0] _T_3654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6918;
  reg [31:0] _T_3654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6919;
  reg [31:0] _T_3655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6920;
  reg [31:0] _T_3655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6921;
  reg [31:0] _T_3656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6922;
  reg [31:0] _T_3656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6923;
  reg [31:0] _T_3657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6924;
  reg [31:0] _T_3657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6925;
  reg [31:0] _T_3658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6926;
  reg [31:0] _T_3658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6927;
  reg [31:0] _T_3659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6928;
  reg [31:0] _T_3659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6929;
  reg [31:0] _T_3660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6930;
  reg [31:0] _T_3660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6931;
  reg [31:0] _T_3661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6932;
  reg [31:0] _T_3661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6933;
  reg [31:0] _T_3662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6934;
  reg [31:0] _T_3662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6935;
  reg [31:0] _T_3663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6936;
  reg [31:0] _T_3663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6937;
  reg [31:0] _T_3664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6938;
  reg [31:0] _T_3664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6939;
  reg [31:0] _T_3665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6940;
  reg [31:0] _T_3665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6941;
  reg [31:0] _T_3666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6942;
  reg [31:0] _T_3666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6943;
  reg [31:0] _T_3667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6944;
  reg [31:0] _T_3667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6945;
  reg [31:0] _T_3668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6946;
  reg [31:0] _T_3668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6947;
  reg [31:0] _T_3669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6948;
  reg [31:0] _T_3669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6949;
  reg [31:0] _T_3670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6950;
  reg [31:0] _T_3670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6951;
  reg [31:0] _T_3671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6952;
  reg [31:0] _T_3671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6953;
  reg [31:0] _T_3672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6954;
  reg [31:0] _T_3672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6955;
  reg [31:0] _T_3673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6956;
  reg [31:0] _T_3673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6957;
  reg [31:0] _T_3674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6958;
  reg [31:0] _T_3674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6959;
  reg [31:0] _T_3675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6960;
  reg [31:0] _T_3675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6961;
  reg [31:0] _T_3676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6962;
  reg [31:0] _T_3676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6963;
  reg [31:0] _T_3677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6964;
  reg [31:0] _T_3677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6965;
  reg [31:0] _T_3678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6966;
  reg [31:0] _T_3678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6967;
  reg [31:0] _T_3679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6968;
  reg [31:0] _T_3679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6969;
  reg [31:0] _T_3680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6970;
  reg [31:0] _T_3680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6971;
  reg [31:0] _T_3681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6972;
  reg [31:0] _T_3681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6973;
  reg [31:0] _T_3682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6974;
  reg [31:0] _T_3682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6975;
  reg [31:0] _T_3683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6976;
  reg [31:0] _T_3683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6977;
  reg [31:0] _T_3684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6978;
  reg [31:0] _T_3684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6979;
  reg [31:0] _T_3685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6980;
  reg [31:0] _T_3685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6981;
  reg [31:0] _T_3686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6982;
  reg [31:0] _T_3686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6983;
  reg [31:0] _T_3687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6984;
  reg [31:0] _T_3687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6985;
  reg [31:0] _T_3688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6986;
  reg [31:0] _T_3688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6987;
  reg [31:0] _T_3689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6988;
  reg [31:0] _T_3689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6989;
  reg [31:0] _T_3690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6990;
  reg [31:0] _T_3690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6991;
  reg [31:0] _T_3691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6992;
  reg [31:0] _T_3691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6993;
  reg [31:0] _T_3692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6994;
  reg [31:0] _T_3692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6995;
  reg [31:0] _T_3693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6996;
  reg [31:0] _T_3693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6997;
  reg [31:0] _T_3694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6998;
  reg [31:0] _T_3694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6999;
  reg [31:0] _T_3695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7000;
  reg [31:0] _T_3695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7001;
  reg [31:0] _T_3696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7002;
  reg [31:0] _T_3696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7003;
  reg [31:0] _T_3697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7004;
  reg [31:0] _T_3697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7005;
  reg [31:0] _T_3698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7006;
  reg [31:0] _T_3698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7007;
  reg [31:0] _T_3699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7008;
  reg [31:0] _T_3699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7009;
  reg [31:0] _T_3700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7010;
  reg [31:0] _T_3700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7011;
  reg [31:0] _T_3701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7012;
  reg [31:0] _T_3701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7013;
  reg [31:0] _T_3702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7014;
  reg [31:0] _T_3702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7015;
  reg [31:0] _T_3703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7016;
  reg [31:0] _T_3703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7017;
  reg [31:0] _T_3704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7018;
  reg [31:0] _T_3704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7019;
  reg [31:0] _T_3705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7020;
  reg [31:0] _T_3705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7021;
  reg [31:0] _T_3706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7022;
  reg [31:0] _T_3706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7023;
  reg [31:0] _T_3707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7024;
  reg [31:0] _T_3707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7025;
  reg [31:0] _T_3708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7026;
  reg [31:0] _T_3708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7027;
  reg [31:0] _T_3709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7028;
  reg [31:0] _T_3709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7029;
  reg [31:0] _T_3710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7030;
  reg [31:0] _T_3710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7031;
  reg [31:0] _T_3711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7032;
  reg [31:0] _T_3711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7033;
  reg [31:0] _T_3712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7034;
  reg [31:0] _T_3712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7035;
  reg [31:0] _T_3713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7036;
  reg [31:0] _T_3713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7037;
  reg [31:0] _T_3714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7038;
  reg [31:0] _T_3714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7039;
  reg [31:0] _T_3715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7040;
  reg [31:0] _T_3715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7041;
  reg [31:0] _T_3716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7042;
  reg [31:0] _T_3716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7043;
  reg [31:0] _T_3717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7044;
  reg [31:0] _T_3717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7045;
  reg [31:0] _T_3718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7046;
  reg [31:0] _T_3718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7047;
  reg [31:0] _T_3719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7048;
  reg [31:0] _T_3719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7049;
  reg [31:0] _T_3720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7050;
  reg [31:0] _T_3720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7051;
  reg [31:0] _T_3721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7052;
  reg [31:0] _T_3721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7053;
  reg [31:0] _T_3722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7054;
  reg [31:0] _T_3722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7055;
  reg [31:0] _T_3723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7056;
  reg [31:0] _T_3723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7057;
  reg [31:0] _T_3724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7058;
  reg [31:0] _T_3724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7059;
  reg [31:0] _T_3725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7060;
  reg [31:0] _T_3725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7061;
  reg [31:0] _T_3726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7062;
  reg [31:0] _T_3726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7063;
  reg [31:0] _T_3727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7064;
  reg [31:0] _T_3727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7065;
  reg [31:0] _T_3728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7066;
  reg [31:0] _T_3728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7067;
  reg [31:0] _T_3729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7068;
  reg [31:0] _T_3729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7069;
  reg [31:0] _T_3730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7070;
  reg [31:0] _T_3730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7071;
  reg [31:0] _T_3731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7072;
  reg [31:0] _T_3731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7073;
  reg [31:0] _T_3732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7074;
  reg [31:0] _T_3732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7075;
  reg [31:0] _T_3733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7076;
  reg [31:0] _T_3733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7077;
  reg [31:0] _T_3734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7078;
  reg [31:0] _T_3734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7079;
  reg [31:0] _T_3735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7080;
  reg [31:0] _T_3735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7081;
  reg [31:0] _T_3736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7082;
  reg [31:0] _T_3736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7083;
  reg [31:0] _T_3737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7084;
  reg [31:0] _T_3737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7085;
  reg [31:0] _T_3738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7086;
  reg [31:0] _T_3738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7087;
  reg [31:0] _T_3739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7088;
  reg [31:0] _T_3739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7089;
  reg [31:0] _T_3740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7090;
  reg [31:0] _T_3740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7091;
  reg [31:0] _T_3741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7092;
  reg [31:0] _T_3741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7093;
  reg [31:0] _T_3742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7094;
  reg [31:0] _T_3742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7095;
  reg [31:0] _T_3743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7096;
  reg [31:0] _T_3743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7097;
  reg [31:0] _T_3744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7098;
  reg [31:0] _T_3744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7099;
  reg [31:0] _T_3745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7100;
  reg [31:0] _T_3745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7101;
  reg [31:0] _T_3746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7102;
  reg [31:0] _T_3746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7103;
  reg [31:0] _T_3747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7104;
  reg [31:0] _T_3747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7105;
  reg [31:0] _T_3748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7106;
  reg [31:0] _T_3748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7107;
  reg [31:0] _T_3749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7108;
  reg [31:0] _T_3749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7109;
  reg [31:0] _T_3750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7110;
  reg [31:0] _T_3750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7111;
  reg [31:0] _T_3751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7112;
  reg [31:0] _T_3751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7113;
  reg [31:0] _T_3752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7114;
  reg [31:0] _T_3752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7115;
  reg [31:0] _T_3753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7116;
  reg [31:0] _T_3753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7117;
  reg [31:0] _T_3754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7118;
  reg [31:0] _T_3754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7119;
  reg [31:0] _T_3755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7120;
  reg [31:0] _T_3755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7121;
  reg [31:0] _T_3756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7122;
  reg [31:0] _T_3756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7123;
  reg [31:0] _T_3757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7124;
  reg [31:0] _T_3757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7125;
  reg [31:0] _T_3758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7126;
  reg [31:0] _T_3758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7127;
  reg [31:0] _T_3759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7128;
  reg [31:0] _T_3759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7129;
  reg [31:0] _T_3760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7130;
  reg [31:0] _T_3760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7131;
  reg [31:0] _T_3761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7132;
  reg [31:0] _T_3761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7133;
  reg [31:0] _T_3762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7134;
  reg [31:0] _T_3762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7135;
  reg [31:0] _T_3763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7136;
  reg [31:0] _T_3763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7137;
  reg [31:0] _T_3764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7138;
  reg [31:0] _T_3764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7139;
  reg [31:0] _T_3765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7140;
  reg [31:0] _T_3765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7141;
  reg [31:0] _T_3766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7142;
  reg [31:0] _T_3766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7143;
  reg [31:0] _T_3767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7144;
  reg [31:0] _T_3767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7145;
  reg [31:0] _T_3768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7146;
  reg [31:0] _T_3768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7147;
  reg [31:0] _T_3769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7148;
  reg [31:0] _T_3769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7149;
  reg [31:0] _T_3770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7150;
  reg [31:0] _T_3770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7151;
  reg [31:0] _T_3771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7152;
  reg [31:0] _T_3771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7153;
  reg [31:0] _T_3772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7154;
  reg [31:0] _T_3772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7155;
  reg [31:0] _T_3773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7156;
  reg [31:0] _T_3773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7157;
  reg [31:0] _T_3774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7158;
  reg [31:0] _T_3774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7159;
  reg [31:0] _T_3775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7160;
  reg [31:0] _T_3775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7161;
  reg [31:0] _T_3776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7162;
  reg [31:0] _T_3776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7163;
  reg [31:0] _T_3777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7164;
  reg [31:0] _T_3777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7165;
  reg [31:0] _T_3778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7166;
  reg [31:0] _T_3778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7167;
  reg [31:0] _T_3779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7168;
  reg [31:0] _T_3779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7169;
  reg [31:0] _T_3780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7170;
  reg [31:0] _T_3780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7171;
  reg [31:0] _T_3781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7172;
  reg [31:0] _T_3781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7173;
  reg [31:0] _T_3782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7174;
  reg [31:0] _T_3782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7175;
  reg [31:0] _T_3783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7176;
  reg [31:0] _T_3783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7177;
  reg [31:0] _T_3784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7178;
  reg [31:0] _T_3784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7179;
  reg [31:0] _T_3785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7180;
  reg [31:0] _T_3785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7181;
  reg [31:0] _T_3786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7182;
  reg [31:0] _T_3786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7183;
  reg [31:0] _T_3787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7184;
  reg [31:0] _T_3787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7185;
  reg [31:0] _T_3788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7186;
  reg [31:0] _T_3788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7187;
  reg [31:0] _T_3789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7188;
  reg [31:0] _T_3789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7189;
  reg [31:0] _T_3790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7190;
  reg [31:0] _T_3790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7191;
  reg [31:0] _T_3791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7192;
  reg [31:0] _T_3791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7193;
  reg [31:0] _T_3792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7194;
  reg [31:0] _T_3792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7195;
  reg [31:0] _T_3793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7196;
  reg [31:0] _T_3793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7197;
  reg [31:0] _T_3794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7198;
  reg [31:0] _T_3794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7199;
  reg [31:0] _T_3795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7200;
  reg [31:0] _T_3795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7201;
  reg [31:0] _T_3796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7202;
  reg [31:0] _T_3796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7203;
  reg [31:0] _T_3797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7204;
  reg [31:0] _T_3797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7205;
  reg [31:0] _T_3798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7206;
  reg [31:0] _T_3798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7207;
  reg [31:0] _T_3799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7208;
  reg [31:0] _T_3799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7209;
  reg [31:0] _T_3800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7210;
  reg [31:0] _T_3800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7211;
  reg [31:0] _T_3801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7212;
  reg [31:0] _T_3801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7213;
  reg [31:0] _T_3802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7214;
  reg [31:0] _T_3802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7215;
  reg [31:0] _T_3803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7216;
  reg [31:0] _T_3803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7217;
  reg [31:0] _T_3804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7218;
  reg [31:0] _T_3804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7219;
  reg [31:0] _T_3805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7220;
  reg [31:0] _T_3805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7221;
  reg [31:0] _T_3806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7222;
  reg [31:0] _T_3806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7223;
  reg [31:0] _T_3807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7224;
  reg [31:0] _T_3807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7225;
  reg [31:0] _T_3808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7226;
  reg [31:0] _T_3808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7227;
  reg [31:0] _T_3809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7228;
  reg [31:0] _T_3809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7229;
  reg [31:0] _T_3810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7230;
  reg [31:0] _T_3810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7231;
  reg [31:0] _T_3811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7232;
  reg [31:0] _T_3811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7233;
  reg [31:0] _T_3812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7234;
  reg [31:0] _T_3812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7235;
  reg [31:0] _T_3813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7236;
  reg [31:0] _T_3813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7237;
  reg [31:0] _T_3814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7238;
  reg [31:0] _T_3814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7239;
  reg [31:0] _T_3815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7240;
  reg [31:0] _T_3815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7241;
  reg [31:0] _T_3816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7242;
  reg [31:0] _T_3816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7243;
  reg [31:0] _T_3817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7244;
  reg [31:0] _T_3817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7245;
  reg [31:0] _T_3818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7246;
  reg [31:0] _T_3818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7247;
  reg [31:0] _T_3819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7248;
  reg [31:0] _T_3819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7249;
  reg [31:0] _T_3820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7250;
  reg [31:0] _T_3820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7251;
  reg [31:0] _T_3821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7252;
  reg [31:0] _T_3821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7253;
  reg [31:0] _T_3822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7254;
  reg [31:0] _T_3822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7255;
  reg [31:0] _T_3823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7256;
  reg [31:0] _T_3823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7257;
  reg [31:0] _T_3824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7258;
  reg [31:0] _T_3824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7259;
  reg [31:0] _T_3825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7260;
  reg [31:0] _T_3825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7261;
  reg [31:0] _T_3826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7262;
  reg [31:0] _T_3826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7263;
  reg [31:0] _T_3827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7264;
  reg [31:0] _T_3827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7265;
  reg [31:0] _T_3828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7266;
  reg [31:0] _T_3828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7267;
  reg [31:0] _T_3829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7268;
  reg [31:0] _T_3829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7269;
  reg [31:0] _T_3830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7270;
  reg [31:0] _T_3830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7271;
  reg [31:0] _T_3831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7272;
  reg [31:0] _T_3831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7273;
  reg [31:0] _T_3832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7274;
  reg [31:0] _T_3832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7275;
  reg [31:0] _T_3833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7276;
  reg [31:0] _T_3833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7277;
  reg [31:0] _T_3834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7278;
  reg [31:0] _T_3834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7279;
  reg [31:0] _T_3835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7280;
  reg [31:0] _T_3835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7281;
  reg [31:0] _T_3836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7282;
  reg [31:0] _T_3836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7283;
  reg [31:0] _T_3837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7284;
  reg [31:0] _T_3837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7285;
  reg [31:0] _T_3838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7286;
  reg [31:0] _T_3838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7287;
  reg [31:0] _T_3839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7288;
  reg [31:0] _T_3839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7289;
  reg [31:0] _T_3840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7290;
  reg [31:0] _T_3840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7291;
  reg [31:0] _T_3841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7292;
  reg [31:0] _T_3841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7293;
  reg [31:0] _T_3842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7294;
  reg [31:0] _T_3842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7295;
  reg [31:0] _T_3843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7296;
  reg [31:0] _T_3843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7297;
  reg [31:0] _T_3844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7298;
  reg [31:0] _T_3844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7299;
  reg [31:0] _T_3845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7300;
  reg [31:0] _T_3845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7301;
  reg [31:0] _T_3846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7302;
  reg [31:0] _T_3846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7303;
  reg [31:0] _T_3847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7304;
  reg [31:0] _T_3847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7305;
  reg [31:0] _T_3848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7306;
  reg [31:0] _T_3848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7307;
  reg [31:0] _T_3849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7308;
  reg [31:0] _T_3849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7309;
  reg [31:0] _T_3850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7310;
  reg [31:0] _T_3850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7311;
  reg [31:0] _T_3851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7312;
  reg [31:0] _T_3851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7313;
  reg [31:0] _T_3852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7314;
  reg [31:0] _T_3852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7315;
  reg [31:0] _T_3853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7316;
  reg [31:0] _T_3853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7317;
  reg [31:0] _T_3854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7318;
  reg [31:0] _T_3854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7319;
  reg [31:0] _T_3855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7320;
  reg [31:0] _T_3855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7321;
  reg [31:0] _T_3856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7322;
  reg [31:0] _T_3856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7323;
  reg [31:0] _T_3857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7324;
  reg [31:0] _T_3857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7325;
  reg [31:0] _T_3858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7326;
  reg [31:0] _T_3858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7327;
  reg [31:0] _T_3859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7328;
  reg [31:0] _T_3859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7329;
  reg [31:0] _T_3860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7330;
  reg [31:0] _T_3860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7331;
  reg [31:0] _T_3861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7332;
  reg [31:0] _T_3861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7333;
  reg [31:0] _T_3862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7334;
  reg [31:0] _T_3862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7335;
  reg [31:0] _T_3863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7336;
  reg [31:0] _T_3863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7337;
  reg [31:0] _T_3864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7338;
  reg [31:0] _T_3864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7339;
  reg [31:0] _T_3865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7340;
  reg [31:0] _T_3865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7341;
  reg [31:0] _T_3866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7342;
  reg [31:0] _T_3866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7343;
  reg [31:0] _T_3867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7344;
  reg [31:0] _T_3867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7345;
  reg [31:0] _T_3868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7346;
  reg [31:0] _T_3868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7347;
  reg [31:0] _T_3869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7348;
  reg [31:0] _T_3869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7349;
  reg [31:0] _T_3870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7350;
  reg [31:0] _T_3870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7351;
  reg [31:0] _T_3871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7352;
  reg [31:0] _T_3871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7353;
  reg [31:0] _T_3872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7354;
  reg [31:0] _T_3872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7355;
  reg [31:0] _T_3873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7356;
  reg [31:0] _T_3873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7357;
  reg [31:0] _T_3874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7358;
  reg [31:0] _T_3874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7359;
  reg [31:0] _T_3875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7360;
  reg [31:0] _T_3875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7361;
  reg [31:0] _T_3876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7362;
  reg [31:0] _T_3876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7363;
  reg [31:0] _T_3877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7364;
  reg [31:0] _T_3877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7365;
  reg [31:0] _T_3878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7366;
  reg [31:0] _T_3878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7367;
  reg [31:0] _T_3879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7368;
  reg [31:0] _T_3879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7369;
  reg [31:0] _T_3880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7370;
  reg [31:0] _T_3880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7371;
  reg [31:0] _T_3881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7372;
  reg [31:0] _T_3881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7373;
  reg [31:0] _T_3882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7374;
  reg [31:0] _T_3882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7375;
  reg [31:0] _T_3883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7376;
  reg [31:0] _T_3883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7377;
  reg [31:0] _T_3884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7378;
  reg [31:0] _T_3884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7379;
  reg [31:0] _T_3885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7380;
  reg [31:0] _T_3885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7381;
  reg [31:0] _T_3886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7382;
  reg [31:0] _T_3886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7383;
  reg [31:0] _T_3887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7384;
  reg [31:0] _T_3887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7385;
  reg [31:0] _T_3888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7386;
  reg [31:0] _T_3888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7387;
  reg [31:0] _T_3889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7388;
  reg [31:0] _T_3889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7389;
  reg [31:0] _T_3890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7390;
  reg [31:0] _T_3890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7391;
  reg [31:0] _T_3891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7392;
  reg [31:0] _T_3891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7393;
  reg [31:0] _T_3892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7394;
  reg [31:0] _T_3892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7395;
  reg [31:0] _T_3893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7396;
  reg [31:0] _T_3893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7397;
  reg [31:0] _T_3894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7398;
  reg [31:0] _T_3894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7399;
  reg [31:0] _T_3895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7400;
  reg [31:0] _T_3895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7401;
  reg [31:0] _T_3896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7402;
  reg [31:0] _T_3896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7403;
  reg [31:0] _T_3897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7404;
  reg [31:0] _T_3897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7405;
  reg [31:0] _T_3898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7406;
  reg [31:0] _T_3898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7407;
  reg [31:0] _T_3899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7408;
  reg [31:0] _T_3899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7409;
  reg [31:0] _T_3900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7410;
  reg [31:0] _T_3900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7411;
  reg [31:0] _T_3901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7412;
  reg [31:0] _T_3901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7413;
  reg [31:0] _T_3902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7414;
  reg [31:0] _T_3902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7415;
  reg [31:0] _T_3903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7416;
  reg [31:0] _T_3903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7417;
  reg [31:0] _T_3904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7418;
  reg [31:0] _T_3904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7419;
  reg [31:0] _T_3905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7420;
  reg [31:0] _T_3905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7421;
  reg [31:0] _T_3906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7422;
  reg [31:0] _T_3906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7423;
  reg [31:0] _T_3907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7424;
  reg [31:0] _T_3907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7425;
  reg [31:0] _T_3908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7426;
  reg [31:0] _T_3908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7427;
  reg [31:0] _T_3909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7428;
  reg [31:0] _T_3909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7429;
  reg [31:0] _T_3910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7430;
  reg [31:0] _T_3910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7431;
  reg [31:0] _T_3911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7432;
  reg [31:0] _T_3911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7433;
  reg [31:0] _T_3912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7434;
  reg [31:0] _T_3912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7435;
  reg [31:0] _T_3913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7436;
  reg [31:0] _T_3913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7437;
  reg [31:0] _T_3914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7438;
  reg [31:0] _T_3914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7439;
  reg [31:0] _T_3915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7440;
  reg [31:0] _T_3915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7441;
  reg [31:0] _T_3916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7442;
  reg [31:0] _T_3916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7443;
  reg [31:0] _T_3917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7444;
  reg [31:0] _T_3917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7445;
  reg [31:0] _T_3918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7446;
  reg [31:0] _T_3918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7447;
  reg [31:0] _T_3919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7448;
  reg [31:0] _T_3919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7449;
  reg [31:0] _T_3920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7450;
  reg [31:0] _T_3920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7451;
  reg [31:0] _T_3921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7452;
  reg [31:0] _T_3921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7453;
  reg [31:0] _T_3922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7454;
  reg [31:0] _T_3922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7455;
  reg [31:0] _T_3923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7456;
  reg [31:0] _T_3923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7457;
  reg [31:0] _T_3924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7458;
  reg [31:0] _T_3924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7459;
  reg [31:0] _T_3925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7460;
  reg [31:0] _T_3925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7461;
  reg [31:0] _T_3926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7462;
  reg [31:0] _T_3926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7463;
  reg [31:0] _T_3927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7464;
  reg [31:0] _T_3927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7465;
  reg [31:0] _T_3928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7466;
  reg [31:0] _T_3928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7467;
  reg [31:0] _T_3929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7468;
  reg [31:0] _T_3929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7469;
  reg [31:0] _T_3930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7470;
  reg [31:0] _T_3930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7471;
  reg [31:0] _T_3931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7472;
  reg [31:0] _T_3931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7473;
  reg [31:0] _T_3932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7474;
  reg [31:0] _T_3932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7475;
  reg [31:0] _T_3933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7476;
  reg [31:0] _T_3933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7477;
  reg [31:0] _T_3934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7478;
  reg [31:0] _T_3934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7479;
  reg [31:0] _T_3935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7480;
  reg [31:0] _T_3935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7481;
  reg [31:0] _T_3936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7482;
  reg [31:0] _T_3936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7483;
  reg [31:0] _T_3937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7484;
  reg [31:0] _T_3937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7485;
  reg [31:0] _T_3938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7486;
  reg [31:0] _T_3938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7487;
  reg [31:0] _T_3939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7488;
  reg [31:0] _T_3939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7489;
  reg [31:0] _T_3940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7490;
  reg [31:0] _T_3940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7491;
  reg [31:0] _T_3941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7492;
  reg [31:0] _T_3941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7493;
  reg [31:0] _T_3942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7494;
  reg [31:0] _T_3942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7495;
  reg [31:0] _T_3943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7496;
  reg [31:0] _T_3943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7497;
  reg [31:0] _T_3944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7498;
  reg [31:0] _T_3944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7499;
  reg [31:0] _T_3945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7500;
  reg [31:0] _T_3945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7501;
  reg [31:0] _T_3946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7502;
  reg [31:0] _T_3946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7503;
  reg [31:0] _T_3947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7504;
  reg [31:0] _T_3947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7505;
  reg [31:0] _T_3948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7506;
  reg [31:0] _T_3948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7507;
  reg [31:0] _T_3949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7508;
  reg [31:0] _T_3949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7509;
  reg [31:0] _T_3950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7510;
  reg [31:0] _T_3950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7511;
  reg [31:0] _T_3951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7512;
  reg [31:0] _T_3951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7513;
  reg [31:0] _T_3952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7514;
  reg [31:0] _T_3952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7515;
  reg [31:0] _T_3953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7516;
  reg [31:0] _T_3953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7517;
  reg [31:0] _T_3954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7518;
  reg [31:0] _T_3954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7519;
  reg [31:0] _T_3955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7520;
  reg [31:0] _T_3955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7521;
  reg [31:0] _T_3956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7522;
  reg [31:0] _T_3956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7523;
  reg [31:0] _T_3957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7524;
  reg [31:0] _T_3957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7525;
  reg [31:0] _T_3958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7526;
  reg [31:0] _T_3958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7527;
  reg [31:0] _T_3959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7528;
  reg [31:0] _T_3959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7529;
  reg [31:0] _T_3960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7530;
  reg [31:0] _T_3960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7531;
  reg [31:0] _T_3961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7532;
  reg [31:0] _T_3961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7533;
  reg [31:0] _T_3962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7534;
  reg [31:0] _T_3962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7535;
  reg [31:0] _T_3963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7536;
  reg [31:0] _T_3963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7537;
  reg [31:0] _T_3964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7538;
  reg [31:0] _T_3964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7539;
  reg [31:0] _T_3965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7540;
  reg [31:0] _T_3965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7541;
  reg [31:0] _T_3966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7542;
  reg [31:0] _T_3966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7543;
  reg [31:0] _T_3967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7544;
  reg [31:0] _T_3967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7545;
  reg [31:0] _T_3968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7546;
  reg [31:0] _T_3968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7547;
  reg [31:0] _T_3969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7548;
  reg [31:0] _T_3969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7549;
  reg [31:0] _T_3970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7550;
  reg [31:0] _T_3970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7551;
  reg [31:0] _T_3971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7552;
  reg [31:0] _T_3971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7553;
  reg [31:0] _T_3972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7554;
  reg [31:0] _T_3972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7555;
  reg [31:0] _T_3973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7556;
  reg [31:0] _T_3973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7557;
  reg [31:0] _T_3974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7558;
  reg [31:0] _T_3974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7559;
  reg [31:0] _T_3975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7560;
  reg [31:0] _T_3975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7561;
  reg [31:0] _T_3976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7562;
  reg [31:0] _T_3976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7563;
  reg [31:0] _T_3977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7564;
  reg [31:0] _T_3977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7565;
  reg [31:0] _T_3978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7566;
  reg [31:0] _T_3978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7567;
  reg [31:0] _T_3979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7568;
  reg [31:0] _T_3979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7569;
  reg [31:0] _T_3980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7570;
  reg [31:0] _T_3980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7571;
  reg [31:0] _T_3981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7572;
  reg [31:0] _T_3981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7573;
  reg [31:0] _T_3982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7574;
  reg [31:0] _T_3982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7575;
  reg [31:0] _T_3983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7576;
  reg [31:0] _T_3983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7577;
  reg [31:0] _T_3984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7578;
  reg [31:0] _T_3984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7579;
  reg [31:0] _T_3985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7580;
  reg [31:0] _T_3985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7581;
  reg [31:0] _T_3986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7582;
  reg [31:0] _T_3986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7583;
  reg [31:0] _T_3987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7584;
  reg [31:0] _T_3987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7585;
  reg [31:0] _T_3988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7586;
  reg [31:0] _T_3988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7587;
  reg [31:0] _T_3989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7588;
  reg [31:0] _T_3989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7589;
  reg [31:0] _T_3990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7590;
  reg [31:0] _T_3990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7591;
  reg [31:0] _T_3991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7592;
  reg [31:0] _T_3991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7593;
  reg [31:0] _T_3992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7594;
  reg [31:0] _T_3992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7595;
  reg [31:0] _T_3993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7596;
  reg [31:0] _T_3993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7597;
  reg [31:0] _T_3994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7598;
  reg [31:0] _T_3994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7599;
  reg [31:0] _T_3995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7600;
  reg [31:0] _T_3995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7601;
  reg [31:0] _T_3996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7602;
  reg [31:0] _T_3996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7603;
  reg [31:0] _T_3997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7604;
  reg [31:0] _T_3997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7605;
  reg [31:0] _T_3998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7606;
  reg [31:0] _T_3998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7607;
  reg [31:0] _T_3999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7608;
  reg [31:0] _T_3999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7609;
  reg [31:0] _T_4000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7610;
  reg [31:0] _T_4000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7611;
  reg [31:0] _T_4001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7612;
  reg [31:0] _T_4001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7613;
  reg [31:0] _T_4002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7614;
  reg [31:0] _T_4002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7615;
  reg [31:0] _T_4003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7616;
  reg [31:0] _T_4003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7617;
  reg [31:0] _T_4004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7618;
  reg [31:0] _T_4004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7619;
  reg [31:0] _T_4005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7620;
  reg [31:0] _T_4005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7621;
  reg [31:0] _T_4006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7622;
  reg [31:0] _T_4006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7623;
  reg [31:0] _T_4007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7624;
  reg [31:0] _T_4007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7625;
  reg [31:0] _T_4008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7626;
  reg [31:0] _T_4008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7627;
  reg [31:0] _T_4009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7628;
  reg [31:0] _T_4009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7629;
  reg [31:0] _T_4010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7630;
  reg [31:0] _T_4010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7631;
  reg [31:0] _T_4011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7632;
  reg [31:0] _T_4011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7633;
  reg [31:0] _T_4012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7634;
  reg [31:0] _T_4012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7635;
  reg [31:0] _T_4013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7636;
  reg [31:0] _T_4013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7637;
  reg [31:0] _T_4014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7638;
  reg [31:0] _T_4014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7639;
  reg [31:0] _T_4015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7640;
  reg [31:0] _T_4015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7641;
  reg [31:0] _T_4016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7642;
  reg [31:0] _T_4016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7643;
  reg [31:0] _T_4017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7644;
  reg [31:0] _T_4017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7645;
  reg [31:0] _T_4018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7646;
  reg [31:0] _T_4018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7647;
  reg [31:0] _T_4019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7648;
  reg [31:0] _T_4019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7649;
  reg [31:0] _T_4020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7650;
  reg [31:0] _T_4020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7651;
  reg [31:0] _T_4021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7652;
  reg [31:0] _T_4021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7653;
  reg [31:0] _T_4022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7654;
  reg [31:0] _T_4022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7655;
  reg [31:0] _T_4023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7656;
  reg [31:0] _T_4023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7657;
  reg [31:0] _T_4024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7658;
  reg [31:0] _T_4024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7659;
  reg [31:0] _T_4025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7660;
  reg [31:0] _T_4025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7661;
  reg [31:0] _T_4026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7662;
  reg [31:0] _T_4026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7663;
  reg [31:0] _T_4027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7664;
  reg [31:0] _T_4027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7665;
  reg [31:0] _T_4028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7666;
  reg [31:0] _T_4028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7667;
  reg [31:0] _T_4029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7668;
  reg [31:0] _T_4029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7669;
  reg [31:0] _T_4030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7670;
  reg [31:0] _T_4030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7671;
  reg [31:0] _T_4031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7672;
  reg [31:0] _T_4031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7673;
  reg [31:0] _T_4032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7674;
  reg [31:0] _T_4032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7675;
  reg [31:0] _T_4033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7676;
  reg [31:0] _T_4033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7677;
  reg [31:0] _T_4034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7678;
  reg [31:0] _T_4034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7679;
  reg [31:0] _T_4035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7680;
  reg [31:0] _T_4035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7681;
  reg [31:0] _T_4036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7682;
  reg [31:0] _T_4036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7683;
  reg [31:0] _T_4037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7684;
  reg [31:0] _T_4037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7685;
  reg [31:0] _T_4038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7686;
  reg [31:0] _T_4038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7687;
  reg [31:0] _T_4039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7688;
  reg [31:0] _T_4039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7689;
  reg [31:0] _T_4040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7690;
  reg [31:0] _T_4040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7691;
  reg [31:0] _T_4041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7692;
  reg [31:0] _T_4041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7693;
  reg [31:0] _T_4042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7694;
  reg [31:0] _T_4042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7695;
  reg [31:0] _T_4043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7696;
  reg [31:0] _T_4043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7697;
  reg [31:0] _T_4044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7698;
  reg [31:0] _T_4044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7699;
  reg [31:0] _T_4045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7700;
  reg [31:0] _T_4045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7701;
  reg [31:0] _T_4046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7702;
  reg [31:0] _T_4046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7703;
  reg [31:0] _T_4047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7704;
  reg [31:0] _T_4047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7705;
  reg [31:0] _T_4048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7706;
  reg [31:0] _T_4048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7707;
  reg [31:0] _T_4049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7708;
  reg [31:0] _T_4049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7709;
  reg [31:0] _T_4050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7710;
  reg [31:0] _T_4050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7711;
  reg [31:0] _T_4051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7712;
  reg [31:0] _T_4051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7713;
  reg [31:0] _T_4052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7714;
  reg [31:0] _T_4052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7715;
  reg [31:0] _T_4053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7716;
  reg [31:0] _T_4053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7717;
  reg [31:0] _T_4054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7718;
  reg [31:0] _T_4054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7719;
  reg [31:0] _T_4055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7720;
  reg [31:0] _T_4055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7721;
  reg [31:0] _T_4056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7722;
  reg [31:0] _T_4056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7723;
  reg [31:0] _T_4057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7724;
  reg [31:0] _T_4057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7725;
  reg [31:0] _T_4058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7726;
  reg [31:0] _T_4058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7727;
  reg [31:0] _T_4059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7728;
  reg [31:0] _T_4059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7729;
  reg [31:0] _T_4060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7730;
  reg [31:0] _T_4060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7731;
  reg [31:0] _T_4061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7732;
  reg [31:0] _T_4061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7733;
  reg [31:0] _T_4062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7734;
  reg [31:0] _T_4062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7735;
  reg [31:0] _T_4063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7736;
  reg [31:0] _T_4063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7737;
  reg [31:0] _T_4064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7738;
  reg [31:0] _T_4064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7739;
  reg [31:0] _T_4065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7740;
  reg [31:0] _T_4065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7741;
  reg [31:0] _T_4066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7742;
  reg [31:0] _T_4066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7743;
  reg [31:0] _T_4067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7744;
  reg [31:0] _T_4067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7745;
  reg [31:0] _T_4068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7746;
  reg [31:0] _T_4068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7747;
  reg [31:0] _T_4069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7748;
  reg [31:0] _T_4069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7749;
  reg [31:0] _T_4070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7750;
  reg [31:0] _T_4070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7751;
  reg [31:0] _T_4071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7752;
  reg [31:0] _T_4071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7753;
  reg [31:0] _T_4072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7754;
  reg [31:0] _T_4072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7755;
  reg [31:0] _T_4073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7756;
  reg [31:0] _T_4073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7757;
  reg [31:0] _T_4074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7758;
  reg [31:0] _T_4074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7759;
  reg [31:0] _T_4075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7760;
  reg [31:0] _T_4075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7761;
  reg [31:0] _T_4076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7762;
  reg [31:0] _T_4076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7763;
  reg [31:0] _T_4077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7764;
  reg [31:0] _T_4077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7765;
  reg [31:0] _T_4078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7766;
  reg [31:0] _T_4078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7767;
  reg [31:0] _T_4079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7768;
  reg [31:0] _T_4079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7769;
  reg [31:0] _T_4080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7770;
  reg [31:0] _T_4080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7771;
  reg [31:0] _T_4081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7772;
  reg [31:0] _T_4081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7773;
  reg [31:0] _T_4082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7774;
  reg [31:0] _T_4082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7775;
  reg [31:0] _T_4083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7776;
  reg [31:0] _T_4083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7777;
  reg [31:0] _T_4084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7778;
  reg [31:0] _T_4084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7779;
  reg [31:0] _T_4085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7780;
  reg [31:0] _T_4085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7781;
  reg [31:0] _T_4086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7782;
  reg [31:0] _T_4086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7783;
  reg [31:0] _T_4087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7784;
  reg [31:0] _T_4087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7785;
  reg [31:0] _T_4088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7786;
  reg [31:0] _T_4088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7787;
  reg [31:0] _T_4089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7788;
  reg [31:0] _T_4089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7789;
  reg [31:0] _T_4090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7790;
  reg [31:0] _T_4090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7791;
  reg [31:0] _T_4091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7792;
  reg [31:0] _T_4091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7793;
  reg [31:0] _T_4092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7794;
  reg [31:0] _T_4092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7795;
  reg [31:0] _T_4093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7796;
  reg [31:0] _T_4093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7797;
  reg [31:0] _T_4094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7798;
  reg [31:0] _T_4094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7799;
  reg [31:0] _T_4095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7800;
  reg [31:0] _T_4095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7801;
  reg [31:0] _T_4096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7802;
  reg [31:0] _T_4096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7803;
  reg [31:0] _T_4097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7804;
  reg [31:0] _T_4097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7805;
  reg [31:0] _T_4098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7806;
  reg [31:0] _T_4098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7807;
  reg [31:0] _T_4099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7808;
  reg [31:0] _T_4099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7809;
  reg [31:0] _T_4100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7810;
  reg [31:0] _T_4100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7811;
  reg [31:0] _T_4101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7812;
  reg [31:0] _T_4101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7813;
  reg [31:0] _T_4102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7814;
  reg [31:0] _T_4102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7815;
  reg [31:0] _T_4103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7816;
  reg [31:0] _T_4103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7817;
  reg [31:0] _T_4104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7818;
  reg [31:0] _T_4104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7819;
  reg [31:0] _T_4105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7820;
  reg [31:0] _T_4105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7821;
  reg [31:0] _T_4106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7822;
  reg [31:0] _T_4106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7823;
  reg [31:0] _T_4107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7824;
  reg [31:0] _T_4107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7825;
  reg [31:0] _T_4108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7826;
  reg [31:0] _T_4108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7827;
  reg [31:0] _T_4109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7828;
  reg [31:0] _T_4109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7829;
  reg [31:0] _T_4110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7830;
  reg [31:0] _T_4110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7831;
  reg [31:0] _T_4111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7832;
  reg [31:0] _T_4111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7833;
  reg [31:0] _T_4112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7834;
  reg [31:0] _T_4112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7835;
  reg [31:0] _T_4113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7836;
  reg [31:0] _T_4113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7837;
  reg [31:0] _T_4114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7838;
  reg [31:0] _T_4114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7839;
  reg [31:0] _T_4115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7840;
  reg [31:0] _T_4115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7841;
  reg [31:0] _T_4116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7842;
  reg [31:0] _T_4116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7843;
  reg [31:0] _T_4117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7844;
  reg [31:0] _T_4117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7845;
  reg [31:0] _T_4118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7846;
  reg [31:0] _T_4118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7847;
  reg [31:0] _T_4119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7848;
  reg [31:0] _T_4119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7849;
  reg [31:0] _T_4120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7850;
  reg [31:0] _T_4120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7851;
  reg [31:0] _T_4121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7852;
  reg [31:0] _T_4121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7853;
  reg [31:0] _T_4122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7854;
  reg [31:0] _T_4122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7855;
  reg [31:0] _T_4123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7856;
  reg [31:0] _T_4123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7857;
  reg [31:0] _T_4124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7858;
  reg [31:0] _T_4124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7859;
  reg [31:0] _T_4125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7860;
  reg [31:0] _T_4125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7861;
  reg [31:0] _T_4126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7862;
  reg [31:0] _T_4126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7863;
  reg [31:0] _T_4127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7864;
  reg [31:0] _T_4127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7865;
  reg [31:0] _T_4128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7866;
  reg [31:0] _T_4128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7867;
  reg [31:0] _T_4129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7868;
  reg [31:0] _T_4129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7869;
  reg [31:0] _T_4130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7870;
  reg [31:0] _T_4130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7871;
  reg [31:0] _T_4131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7872;
  reg [31:0] _T_4131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7873;
  reg [31:0] _T_4132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7874;
  reg [31:0] _T_4132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7875;
  reg [31:0] _T_4133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7876;
  reg [31:0] _T_4133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7877;
  reg [31:0] _T_4134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7878;
  reg [31:0] _T_4134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7879;
  reg [31:0] _T_4135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7880;
  reg [31:0] _T_4135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7881;
  reg [31:0] _T_4136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7882;
  reg [31:0] _T_4136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7883;
  reg [31:0] _T_4137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7884;
  reg [31:0] _T_4137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7885;
  reg [31:0] _T_4138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7886;
  reg [31:0] _T_4138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7887;
  reg [31:0] _T_4139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7888;
  reg [31:0] _T_4139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7889;
  reg [31:0] _T_4140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7890;
  reg [31:0] _T_4140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7891;
  reg [31:0] _T_4141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7892;
  reg [31:0] _T_4141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7893;
  reg [31:0] _T_4142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7894;
  reg [31:0] _T_4142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7895;
  reg [31:0] _T_4143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7896;
  reg [31:0] _T_4143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7897;
  reg [31:0] _T_4144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7898;
  reg [31:0] _T_4144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7899;
  reg [31:0] _T_4145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7900;
  reg [31:0] _T_4145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7901;
  reg [31:0] _T_4146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7902;
  reg [31:0] _T_4146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7903;
  reg [31:0] _T_4147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7904;
  reg [31:0] _T_4147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7905;
  reg [31:0] _T_4148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7906;
  reg [31:0] _T_4148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7907;
  reg [31:0] _T_4149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7908;
  reg [31:0] _T_4149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7909;
  reg [31:0] _T_4150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7910;
  reg [31:0] _T_4150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7911;
  reg [31:0] _T_4151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7912;
  reg [31:0] _T_4151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7913;
  reg [31:0] _T_4152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7914;
  reg [31:0] _T_4152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7915;
  reg [31:0] _T_4153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7916;
  reg [31:0] _T_4153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7917;
  reg [31:0] _T_4154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7918;
  reg [31:0] _T_4154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7919;
  reg [31:0] _T_4155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7920;
  reg [31:0] _T_4155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7921;
  reg [31:0] _T_4156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7922;
  reg [31:0] _T_4156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7923;
  reg [31:0] _T_4157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7924;
  reg [31:0] _T_4157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7925;
  reg [31:0] _T_4158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7926;
  reg [31:0] _T_4158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7927;
  reg [31:0] _T_4159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7928;
  reg [31:0] _T_4159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7929;
  reg [31:0] _T_4160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7930;
  reg [31:0] _T_4160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7931;
  reg [31:0] _T_4161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7932;
  reg [31:0] _T_4161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7933;
  reg [31:0] _T_4162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7934;
  reg [31:0] _T_4162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7935;
  reg [31:0] _T_4163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7936;
  reg [31:0] _T_4163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7937;
  reg [31:0] _T_4164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7938;
  reg [31:0] _T_4164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7939;
  reg [31:0] _T_4165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7940;
  reg [31:0] _T_4165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7941;
  reg [31:0] _T_4166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7942;
  reg [31:0] _T_4166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7943;
  reg [31:0] _T_4167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7944;
  reg [31:0] _T_4167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7945;
  reg [31:0] _T_4168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7946;
  reg [31:0] _T_4168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7947;
  reg [31:0] _T_4169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7948;
  reg [31:0] _T_4169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7949;
  reg [31:0] _T_4170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7950;
  reg [31:0] _T_4170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7951;
  reg [31:0] _T_4171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7952;
  reg [31:0] _T_4171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7953;
  reg [31:0] _T_4172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7954;
  reg [31:0] _T_4172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7955;
  reg [31:0] _T_4173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7956;
  reg [31:0] _T_4173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7957;
  reg [31:0] _T_4174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7958;
  reg [31:0] _T_4174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7959;
  reg [31:0] _T_4175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7960;
  reg [31:0] _T_4175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7961;
  reg [31:0] _T_4176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7962;
  reg [31:0] _T_4176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7963;
  reg [31:0] _T_4177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7964;
  reg [31:0] _T_4177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7965;
  reg [31:0] _T_4178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7966;
  reg [31:0] _T_4178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7967;
  reg [31:0] _T_4179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7968;
  reg [31:0] _T_4179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7969;
  reg [31:0] _T_4180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7970;
  reg [31:0] _T_4180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7971;
  reg [31:0] _T_4181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7972;
  reg [31:0] _T_4181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7973;
  reg [31:0] _T_4182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7974;
  reg [31:0] _T_4182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7975;
  reg [31:0] _T_4183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7976;
  reg [31:0] _T_4183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7977;
  reg [31:0] _T_4184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7978;
  reg [31:0] _T_4184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7979;
  reg [31:0] _T_4185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7980;
  reg [31:0] _T_4185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7981;
  reg [31:0] _T_4186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7982;
  reg [31:0] _T_4186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7983;
  reg [31:0] _T_4187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7984;
  reg [31:0] _T_4187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7985;
  reg [31:0] _T_4188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7986;
  reg [31:0] _T_4188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7987;
  reg [31:0] _T_4189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7988;
  reg [31:0] _T_4189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7989;
  reg [31:0] _T_4190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7990;
  reg [31:0] _T_4190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7991;
  reg [31:0] _T_4191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7992;
  reg [31:0] _T_4191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7993;
  reg [31:0] _T_4192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7994;
  reg [31:0] _T_4192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7995;
  reg [31:0] _T_4193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7996;
  reg [31:0] _T_4193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7997;
  reg [31:0] _T_4194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7998;
  reg [31:0] _T_4194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7999;
  reg [31:0] _T_4195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8000;
  reg [31:0] _T_4195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8001;
  reg [31:0] _T_4196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8002;
  reg [31:0] _T_4196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8003;
  reg [31:0] _T_4197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8004;
  reg [31:0] _T_4197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8005;
  reg [31:0] _T_4198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8006;
  reg [31:0] _T_4198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8007;
  reg [31:0] _T_4199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8008;
  reg [31:0] _T_4199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8009;
  reg [31:0] _T_4200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8010;
  reg [31:0] _T_4200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8011;
  reg [31:0] _T_4201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8012;
  reg [31:0] _T_4201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8013;
  reg [31:0] _T_4202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8014;
  reg [31:0] _T_4202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8015;
  reg [31:0] _T_4203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8016;
  reg [31:0] _T_4203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8017;
  reg [31:0] _T_4204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8018;
  reg [31:0] _T_4204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8019;
  reg [31:0] _T_4205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8020;
  reg [31:0] _T_4205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8021;
  reg [31:0] _T_4206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8022;
  reg [31:0] _T_4206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8023;
  reg [31:0] _T_4207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8024;
  reg [31:0] _T_4207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8025;
  reg [31:0] _T_4208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8026;
  reg [31:0] _T_4208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8027;
  reg [31:0] _T_4209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8028;
  reg [31:0] _T_4209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8029;
  reg [31:0] _T_4210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8030;
  reg [31:0] _T_4210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8031;
  reg [31:0] _T_4211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8032;
  reg [31:0] _T_4211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8033;
  reg [31:0] _T_4212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8034;
  reg [31:0] _T_4212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8035;
  reg [31:0] _T_4213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8036;
  reg [31:0] _T_4213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8037;
  reg [31:0] _T_4214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8038;
  reg [31:0] _T_4214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8039;
  reg [31:0] _T_4215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8040;
  reg [31:0] _T_4215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8041;
  reg [31:0] _T_4216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8042;
  reg [31:0] _T_4216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8043;
  reg [31:0] _T_4217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8044;
  reg [31:0] _T_4217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8045;
  reg [31:0] _T_4218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8046;
  reg [31:0] _T_4218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8047;
  reg [31:0] _T_4219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8048;
  reg [31:0] _T_4219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8049;
  reg [31:0] _T_4220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8050;
  reg [31:0] _T_4220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8051;
  reg [31:0] _T_4221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8052;
  reg [31:0] _T_4221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8053;
  reg [31:0] _T_4222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8054;
  reg [31:0] _T_4222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8055;
  reg [31:0] _T_4223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8056;
  reg [31:0] _T_4223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8057;
  reg [31:0] _T_4224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8058;
  reg [31:0] _T_4224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8059;
  reg [31:0] _T_4225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8060;
  reg [31:0] _T_4225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8061;
  reg [31:0] _T_4226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8062;
  reg [31:0] _T_4226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8063;
  reg [31:0] _T_4227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8064;
  reg [31:0] _T_4227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8065;
  reg [31:0] _T_4228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8066;
  reg [31:0] _T_4228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8067;
  reg [31:0] _T_4229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8068;
  reg [31:0] _T_4229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8069;
  reg [31:0] _T_4230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8070;
  reg [31:0] _T_4230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8071;
  reg [31:0] _T_4231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8072;
  reg [31:0] _T_4231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8073;
  reg [31:0] _T_4232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8074;
  reg [31:0] _T_4232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8075;
  reg [31:0] _T_4233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8076;
  reg [31:0] _T_4233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8077;
  reg [31:0] _T_4234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8078;
  reg [31:0] _T_4234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8079;
  reg [31:0] _T_4235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8080;
  reg [31:0] _T_4235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8081;
  reg [31:0] _T_4236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8082;
  reg [31:0] _T_4236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8083;
  reg [31:0] _T_4237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8084;
  reg [31:0] _T_4237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8085;
  reg [31:0] _T_4238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8086;
  reg [31:0] _T_4238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8087;
  reg [31:0] _T_4239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8088;
  reg [31:0] _T_4239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8089;
  reg [31:0] _T_4240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8090;
  reg [31:0] _T_4240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8091;
  reg [31:0] _T_4241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8092;
  reg [31:0] _T_4241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8093;
  reg [31:0] _T_4242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8094;
  reg [31:0] _T_4242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8095;
  reg [31:0] _T_4243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8096;
  reg [31:0] _T_4243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8097;
  reg [31:0] _T_4244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8098;
  reg [31:0] _T_4244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8099;
  reg [31:0] _T_4245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8100;
  reg [31:0] _T_4245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8101;
  reg [31:0] _T_4246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8102;
  reg [31:0] _T_4246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8103;
  reg [31:0] _T_4247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8104;
  reg [31:0] _T_4247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8105;
  reg [31:0] _T_4248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8106;
  reg [31:0] _T_4248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8107;
  reg [31:0] _T_4249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8108;
  reg [31:0] _T_4249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8109;
  reg [31:0] _T_4250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8110;
  reg [31:0] _T_4250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8111;
  reg [31:0] _T_4251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8112;
  reg [31:0] _T_4251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8113;
  reg [31:0] _T_4252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8114;
  reg [31:0] _T_4252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8115;
  reg [31:0] _T_4253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8116;
  reg [31:0] _T_4253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8117;
  reg [31:0] _T_4254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8118;
  reg [31:0] _T_4254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8119;
  reg [31:0] _T_4255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8120;
  reg [31:0] _T_4255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8121;
  reg [31:0] _T_4256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8122;
  reg [31:0] _T_4256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8123;
  reg [31:0] _T_4257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8124;
  reg [31:0] _T_4257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8125;
  reg [31:0] _T_4258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8126;
  reg [31:0] _T_4258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8127;
  reg [31:0] _T_4259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8128;
  reg [31:0] _T_4259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8129;
  reg [31:0] _T_4260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8130;
  reg [31:0] _T_4260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8131;
  reg [31:0] _T_4261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8132;
  reg [31:0] _T_4261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8133;
  reg [31:0] _T_4262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8134;
  reg [31:0] _T_4262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8135;
  reg [31:0] _T_4263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8136;
  reg [31:0] _T_4263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8137;
  reg [31:0] _T_4264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8138;
  reg [31:0] _T_4264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8139;
  reg [31:0] _T_4265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8140;
  reg [31:0] _T_4265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8141;
  reg [31:0] _T_4266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8142;
  reg [31:0] _T_4266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8143;
  reg [31:0] _T_4267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8144;
  reg [31:0] _T_4267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8145;
  reg [31:0] _T_4268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8146;
  reg [31:0] _T_4268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8147;
  reg [31:0] _T_4269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8148;
  reg [31:0] _T_4269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8149;
  reg [31:0] _T_4270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8150;
  reg [31:0] _T_4270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8151;
  reg [31:0] _T_4271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8152;
  reg [31:0] _T_4271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8153;
  reg [31:0] _T_4272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8154;
  reg [31:0] _T_4272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8155;
  reg [31:0] _T_4273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8156;
  reg [31:0] _T_4273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8157;
  reg [31:0] _T_4274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8158;
  reg [31:0] _T_4274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8159;
  reg [31:0] _T_4275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8160;
  reg [31:0] _T_4275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8161;
  reg [31:0] _T_4276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8162;
  reg [31:0] _T_4276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8163;
  reg [31:0] _T_4277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8164;
  reg [31:0] _T_4277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8165;
  reg [31:0] _T_4278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8166;
  reg [31:0] _T_4278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8167;
  reg [31:0] _T_4279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8168;
  reg [31:0] _T_4279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8169;
  reg [31:0] _T_4280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8170;
  reg [31:0] _T_4280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8171;
  reg [31:0] _T_4281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8172;
  reg [31:0] _T_4281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8173;
  reg [31:0] _T_4282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8174;
  reg [31:0] _T_4282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8175;
  reg [31:0] _T_4283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8176;
  reg [31:0] _T_4283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8177;
  reg [31:0] _T_4284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8178;
  reg [31:0] _T_4284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8179;
  reg [31:0] _T_4285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8180;
  reg [31:0] _T_4285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8181;
  reg [31:0] _T_4286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8182;
  reg [31:0] _T_4286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8183;
  reg [31:0] _T_4287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8184;
  reg [31:0] _T_4287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8185;
  reg [31:0] _T_4288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8186;
  reg [31:0] _T_4288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8187;
  reg [31:0] _T_4289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8188;
  reg [31:0] _T_4289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8189;
  reg [31:0] _T_4290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8190;
  reg [31:0] _T_4290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8191;
  reg [31:0] _T_4291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8192;
  reg [31:0] _T_4291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8193;
  reg [31:0] _T_4294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8194;
  reg [31:0] _T_4294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8195;
  reg [31:0] _T_4295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8196;
  reg [31:0] _T_4295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8197;
  reg [31:0] _T_4296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8198;
  reg [31:0] _T_4296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8199;
  reg [31:0] _T_4297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8200;
  reg [31:0] _T_4297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8201;
  reg [31:0] _T_4298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8202;
  reg [31:0] _T_4298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8203;
  reg [31:0] _T_4299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8204;
  reg [31:0] _T_4299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8205;
  reg [31:0] _T_4300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8206;
  reg [31:0] _T_4300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8207;
  reg [31:0] _T_4301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8208;
  reg [31:0] _T_4301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8209;
  reg [31:0] _T_4302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8210;
  reg [31:0] _T_4302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8211;
  reg [31:0] _T_4303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8212;
  reg [31:0] _T_4303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8213;
  reg [31:0] _T_4304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8214;
  reg [31:0] _T_4304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8215;
  reg [31:0] _T_4305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8216;
  reg [31:0] _T_4305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8217;
  reg [31:0] _T_4306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8218;
  reg [31:0] _T_4306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8219;
  reg [31:0] _T_4307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8220;
  reg [31:0] _T_4307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8221;
  reg [31:0] _T_4308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8222;
  reg [31:0] _T_4308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8223;
  reg [31:0] _T_4309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8224;
  reg [31:0] _T_4309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8225;
  reg [31:0] _T_4310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8226;
  reg [31:0] _T_4310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8227;
  reg [31:0] _T_4311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8228;
  reg [31:0] _T_4311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8229;
  reg [31:0] _T_4312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8230;
  reg [31:0] _T_4312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8231;
  reg [31:0] _T_4313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8232;
  reg [31:0] _T_4313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8233;
  reg [31:0] _T_4314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8234;
  reg [31:0] _T_4314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8235;
  reg [31:0] _T_4315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8236;
  reg [31:0] _T_4315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8237;
  reg [31:0] _T_4316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8238;
  reg [31:0] _T_4316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8239;
  reg [31:0] _T_4317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8240;
  reg [31:0] _T_4317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8241;
  reg [31:0] _T_4318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8242;
  reg [31:0] _T_4318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8243;
  reg [31:0] _T_4319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8244;
  reg [31:0] _T_4319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8245;
  reg [31:0] _T_4320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8246;
  reg [31:0] _T_4320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8247;
  reg [31:0] _T_4321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8248;
  reg [31:0] _T_4321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8249;
  reg [31:0] _T_4322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8250;
  reg [31:0] _T_4322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8251;
  reg [31:0] _T_4323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8252;
  reg [31:0] _T_4323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8253;
  reg [31:0] _T_4324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8254;
  reg [31:0] _T_4324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8255;
  reg [31:0] _T_4325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8256;
  reg [31:0] _T_4325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8257;
  reg [31:0] _T_4326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8258;
  reg [31:0] _T_4326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8259;
  reg [31:0] _T_4327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8260;
  reg [31:0] _T_4327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8261;
  reg [31:0] _T_4328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8262;
  reg [31:0] _T_4328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8263;
  reg [31:0] _T_4329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8264;
  reg [31:0] _T_4329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8265;
  reg [31:0] _T_4330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8266;
  reg [31:0] _T_4330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8267;
  reg [31:0] _T_4331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8268;
  reg [31:0] _T_4331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8269;
  reg [31:0] _T_4332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8270;
  reg [31:0] _T_4332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8271;
  reg [31:0] _T_4333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8272;
  reg [31:0] _T_4333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8273;
  reg [31:0] _T_4334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8274;
  reg [31:0] _T_4334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8275;
  reg [31:0] _T_4335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8276;
  reg [31:0] _T_4335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8277;
  reg [31:0] _T_4336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8278;
  reg [31:0] _T_4336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8279;
  reg [31:0] _T_4337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8280;
  reg [31:0] _T_4337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8281;
  reg [31:0] _T_4338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8282;
  reg [31:0] _T_4338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8283;
  reg [31:0] _T_4339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8284;
  reg [31:0] _T_4339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8285;
  reg [31:0] _T_4340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8286;
  reg [31:0] _T_4340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8287;
  reg [31:0] _T_4341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8288;
  reg [31:0] _T_4341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8289;
  reg [31:0] _T_4342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8290;
  reg [31:0] _T_4342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8291;
  reg [31:0] _T_4343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8292;
  reg [31:0] _T_4343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8293;
  reg [31:0] _T_4344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8294;
  reg [31:0] _T_4344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8295;
  reg [31:0] _T_4345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8296;
  reg [31:0] _T_4345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8297;
  reg [31:0] _T_4346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8298;
  reg [31:0] _T_4346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8299;
  reg [31:0] _T_4347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8300;
  reg [31:0] _T_4347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8301;
  reg [31:0] _T_4348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8302;
  reg [31:0] _T_4348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8303;
  reg [31:0] _T_4349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8304;
  reg [31:0] _T_4349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8305;
  reg [31:0] _T_4350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8306;
  reg [31:0] _T_4350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8307;
  reg [31:0] _T_4351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8308;
  reg [31:0] _T_4351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8309;
  reg [31:0] _T_4352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8310;
  reg [31:0] _T_4352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8311;
  reg [31:0] _T_4353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8312;
  reg [31:0] _T_4353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8313;
  reg [31:0] _T_4354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8314;
  reg [31:0] _T_4354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8315;
  reg [31:0] _T_4355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8316;
  reg [31:0] _T_4355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8317;
  reg [31:0] _T_4356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8318;
  reg [31:0] _T_4356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8319;
  reg [31:0] _T_4357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8320;
  reg [31:0] _T_4357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8321;
  reg [31:0] _T_4358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8322;
  reg [31:0] _T_4358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8323;
  reg [31:0] _T_4359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8324;
  reg [31:0] _T_4359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8325;
  reg [31:0] _T_4360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8326;
  reg [31:0] _T_4360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8327;
  reg [31:0] _T_4361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8328;
  reg [31:0] _T_4361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8329;
  reg [31:0] _T_4362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8330;
  reg [31:0] _T_4362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8331;
  reg [31:0] _T_4363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8332;
  reg [31:0] _T_4363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8333;
  reg [31:0] _T_4364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8334;
  reg [31:0] _T_4364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8335;
  reg [31:0] _T_4365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8336;
  reg [31:0] _T_4365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8337;
  reg [31:0] _T_4366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8338;
  reg [31:0] _T_4366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8339;
  reg [31:0] _T_4367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8340;
  reg [31:0] _T_4367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8341;
  reg [31:0] _T_4368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8342;
  reg [31:0] _T_4368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8343;
  reg [31:0] _T_4369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8344;
  reg [31:0] _T_4369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8345;
  reg [31:0] _T_4370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8346;
  reg [31:0] _T_4370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8347;
  reg [31:0] _T_4371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8348;
  reg [31:0] _T_4371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8349;
  reg [31:0] _T_4372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8350;
  reg [31:0] _T_4372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8351;
  reg [31:0] _T_4373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8352;
  reg [31:0] _T_4373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8353;
  reg [31:0] _T_4374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8354;
  reg [31:0] _T_4374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8355;
  reg [31:0] _T_4375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8356;
  reg [31:0] _T_4375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8357;
  reg [31:0] _T_4376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8358;
  reg [31:0] _T_4376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8359;
  reg [31:0] _T_4377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8360;
  reg [31:0] _T_4377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8361;
  reg [31:0] _T_4378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8362;
  reg [31:0] _T_4378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8363;
  reg [31:0] _T_4379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8364;
  reg [31:0] _T_4379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8365;
  reg [31:0] _T_4380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8366;
  reg [31:0] _T_4380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8367;
  reg [31:0] _T_4381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8368;
  reg [31:0] _T_4381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8369;
  reg [31:0] _T_4382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8370;
  reg [31:0] _T_4382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8371;
  reg [31:0] _T_4383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8372;
  reg [31:0] _T_4383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8373;
  reg [31:0] _T_4384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8374;
  reg [31:0] _T_4384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8375;
  reg [31:0] _T_4385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8376;
  reg [31:0] _T_4385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8377;
  reg [31:0] _T_4386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8378;
  reg [31:0] _T_4386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8379;
  reg [31:0] _T_4387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8380;
  reg [31:0] _T_4387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8381;
  reg [31:0] _T_4388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8382;
  reg [31:0] _T_4388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8383;
  reg [31:0] _T_4389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8384;
  reg [31:0] _T_4389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8385;
  reg [31:0] _T_4390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8386;
  reg [31:0] _T_4390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8387;
  reg [31:0] _T_4391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8388;
  reg [31:0] _T_4391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8389;
  reg [31:0] _T_4392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8390;
  reg [31:0] _T_4392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8391;
  reg [31:0] _T_4393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8392;
  reg [31:0] _T_4393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8393;
  reg [31:0] _T_4394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8394;
  reg [31:0] _T_4394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8395;
  reg [31:0] _T_4395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8396;
  reg [31:0] _T_4395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8397;
  reg [31:0] _T_4396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8398;
  reg [31:0] _T_4396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8399;
  reg [31:0] _T_4397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8400;
  reg [31:0] _T_4397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8401;
  reg [31:0] _T_4398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8402;
  reg [31:0] _T_4398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8403;
  reg [31:0] _T_4399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8404;
  reg [31:0] _T_4399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8405;
  reg [31:0] _T_4400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8406;
  reg [31:0] _T_4400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8407;
  reg [31:0] _T_4401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8408;
  reg [31:0] _T_4401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8409;
  reg [31:0] _T_4402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8410;
  reg [31:0] _T_4402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8411;
  reg [31:0] _T_4403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8412;
  reg [31:0] _T_4403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8413;
  reg [31:0] _T_4404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8414;
  reg [31:0] _T_4404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8415;
  reg [31:0] _T_4405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8416;
  reg [31:0] _T_4405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8417;
  reg [31:0] _T_4406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8418;
  reg [31:0] _T_4406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8419;
  reg [31:0] _T_4407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8420;
  reg [31:0] _T_4407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8421;
  reg [31:0] _T_4408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8422;
  reg [31:0] _T_4408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8423;
  reg [31:0] _T_4409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8424;
  reg [31:0] _T_4409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8425;
  reg [31:0] _T_4410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8426;
  reg [31:0] _T_4410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8427;
  reg [31:0] _T_4411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8428;
  reg [31:0] _T_4411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8429;
  reg [31:0] _T_4412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8430;
  reg [31:0] _T_4412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8431;
  reg [31:0] _T_4413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8432;
  reg [31:0] _T_4413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8433;
  reg [31:0] _T_4414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8434;
  reg [31:0] _T_4414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8435;
  reg [31:0] _T_4415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8436;
  reg [31:0] _T_4415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8437;
  reg [31:0] _T_4416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8438;
  reg [31:0] _T_4416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8439;
  reg [31:0] _T_4417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8440;
  reg [31:0] _T_4417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8441;
  reg [31:0] _T_4418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8442;
  reg [31:0] _T_4418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8443;
  reg [31:0] _T_4419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8444;
  reg [31:0] _T_4419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8445;
  reg [31:0] _T_4420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8446;
  reg [31:0] _T_4420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8447;
  reg [31:0] _T_4421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8448;
  reg [31:0] _T_4421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8449;
  reg [31:0] _T_4422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8450;
  reg [31:0] _T_4422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8451;
  reg [31:0] _T_4423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8452;
  reg [31:0] _T_4423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8453;
  reg [31:0] _T_4424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8454;
  reg [31:0] _T_4424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8455;
  reg [31:0] _T_4425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8456;
  reg [31:0] _T_4425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8457;
  reg [31:0] _T_4426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8458;
  reg [31:0] _T_4426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8459;
  reg [31:0] _T_4427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8460;
  reg [31:0] _T_4427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8461;
  reg [31:0] _T_4428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8462;
  reg [31:0] _T_4428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8463;
  reg [31:0] _T_4429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8464;
  reg [31:0] _T_4429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8465;
  reg [31:0] _T_4430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8466;
  reg [31:0] _T_4430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8467;
  reg [31:0] _T_4431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8468;
  reg [31:0] _T_4431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8469;
  reg [31:0] _T_4432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8470;
  reg [31:0] _T_4432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8471;
  reg [31:0] _T_4433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8472;
  reg [31:0] _T_4433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8473;
  reg [31:0] _T_4434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8474;
  reg [31:0] _T_4434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8475;
  reg [31:0] _T_4435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8476;
  reg [31:0] _T_4435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8477;
  reg [31:0] _T_4436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8478;
  reg [31:0] _T_4436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8479;
  reg [31:0] _T_4437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8480;
  reg [31:0] _T_4437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8481;
  reg [31:0] _T_4438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8482;
  reg [31:0] _T_4438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8483;
  reg [31:0] _T_4439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8484;
  reg [31:0] _T_4439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8485;
  reg [31:0] _T_4440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8486;
  reg [31:0] _T_4440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8487;
  reg [31:0] _T_4441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8488;
  reg [31:0] _T_4441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8489;
  reg [31:0] _T_4442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8490;
  reg [31:0] _T_4442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8491;
  reg [31:0] _T_4443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8492;
  reg [31:0] _T_4443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8493;
  reg [31:0] _T_4444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8494;
  reg [31:0] _T_4444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8495;
  reg [31:0] _T_4445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8496;
  reg [31:0] _T_4445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8497;
  reg [31:0] _T_4446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8498;
  reg [31:0] _T_4446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8499;
  reg [31:0] _T_4447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8500;
  reg [31:0] _T_4447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8501;
  reg [31:0] _T_4448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8502;
  reg [31:0] _T_4448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8503;
  reg [31:0] _T_4449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8504;
  reg [31:0] _T_4449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8505;
  reg [31:0] _T_4450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8506;
  reg [31:0] _T_4450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8507;
  reg [31:0] _T_4451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8508;
  reg [31:0] _T_4451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8509;
  reg [31:0] _T_4452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8510;
  reg [31:0] _T_4452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8511;
  reg [31:0] _T_4453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8512;
  reg [31:0] _T_4453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8513;
  reg [31:0] _T_4454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8514;
  reg [31:0] _T_4454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8515;
  reg [31:0] _T_4455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8516;
  reg [31:0] _T_4455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8517;
  reg [31:0] _T_4456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8518;
  reg [31:0] _T_4456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8519;
  reg [31:0] _T_4457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8520;
  reg [31:0] _T_4457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8521;
  reg [31:0] _T_4458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8522;
  reg [31:0] _T_4458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8523;
  reg [31:0] _T_4459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8524;
  reg [31:0] _T_4459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8525;
  reg [31:0] _T_4460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8526;
  reg [31:0] _T_4460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8527;
  reg [31:0] _T_4461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8528;
  reg [31:0] _T_4461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8529;
  reg [31:0] _T_4462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8530;
  reg [31:0] _T_4462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8531;
  reg [31:0] _T_4463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8532;
  reg [31:0] _T_4463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8533;
  reg [31:0] _T_4464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8534;
  reg [31:0] _T_4464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8535;
  reg [31:0] _T_4465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8536;
  reg [31:0] _T_4465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8537;
  reg [31:0] _T_4466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8538;
  reg [31:0] _T_4466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8539;
  reg [31:0] _T_4467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8540;
  reg [31:0] _T_4467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8541;
  reg [31:0] _T_4468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8542;
  reg [31:0] _T_4468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8543;
  reg [31:0] _T_4469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8544;
  reg [31:0] _T_4469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8545;
  reg [31:0] _T_4470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8546;
  reg [31:0] _T_4470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8547;
  reg [31:0] _T_4471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8548;
  reg [31:0] _T_4471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8549;
  reg [31:0] _T_4472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8550;
  reg [31:0] _T_4472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8551;
  reg [31:0] _T_4473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8552;
  reg [31:0] _T_4473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8553;
  reg [31:0] _T_4474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8554;
  reg [31:0] _T_4474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8555;
  reg [31:0] _T_4475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8556;
  reg [31:0] _T_4475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8557;
  reg [31:0] _T_4476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8558;
  reg [31:0] _T_4476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8559;
  reg [31:0] _T_4477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8560;
  reg [31:0] _T_4477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8561;
  reg [31:0] _T_4478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8562;
  reg [31:0] _T_4478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8563;
  reg [31:0] _T_4479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8564;
  reg [31:0] _T_4479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8565;
  reg [31:0] _T_4480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8566;
  reg [31:0] _T_4480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8567;
  reg [31:0] _T_4481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8568;
  reg [31:0] _T_4481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8569;
  reg [31:0] _T_4482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8570;
  reg [31:0] _T_4482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8571;
  reg [31:0] _T_4483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8572;
  reg [31:0] _T_4483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8573;
  reg [31:0] _T_4484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8574;
  reg [31:0] _T_4484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8575;
  reg [31:0] _T_4485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8576;
  reg [31:0] _T_4485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8577;
  reg [31:0] _T_4486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8578;
  reg [31:0] _T_4486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8579;
  reg [31:0] _T_4487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8580;
  reg [31:0] _T_4487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8581;
  reg [31:0] _T_4488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8582;
  reg [31:0] _T_4488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8583;
  reg [31:0] _T_4489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8584;
  reg [31:0] _T_4489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8585;
  reg [31:0] _T_4490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8586;
  reg [31:0] _T_4490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8587;
  reg [31:0] _T_4491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8588;
  reg [31:0] _T_4491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8589;
  reg [31:0] _T_4492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8590;
  reg [31:0] _T_4492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8591;
  reg [31:0] _T_4493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8592;
  reg [31:0] _T_4493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8593;
  reg [31:0] _T_4494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8594;
  reg [31:0] _T_4494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8595;
  reg [31:0] _T_4495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8596;
  reg [31:0] _T_4495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8597;
  reg [31:0] _T_4496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8598;
  reg [31:0] _T_4496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8599;
  reg [31:0] _T_4497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8600;
  reg [31:0] _T_4497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8601;
  reg [31:0] _T_4498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8602;
  reg [31:0] _T_4498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8603;
  reg [31:0] _T_4499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8604;
  reg [31:0] _T_4499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8605;
  reg [31:0] _T_4500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8606;
  reg [31:0] _T_4500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8607;
  reg [31:0] _T_4501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8608;
  reg [31:0] _T_4501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8609;
  reg [31:0] _T_4502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8610;
  reg [31:0] _T_4502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8611;
  reg [31:0] _T_4503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8612;
  reg [31:0] _T_4503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8613;
  reg [31:0] _T_4504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8614;
  reg [31:0] _T_4504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8615;
  reg [31:0] _T_4505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8616;
  reg [31:0] _T_4505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8617;
  reg [31:0] _T_4506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8618;
  reg [31:0] _T_4506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8619;
  reg [31:0] _T_4507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8620;
  reg [31:0] _T_4507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8621;
  reg [31:0] _T_4508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8622;
  reg [31:0] _T_4508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8623;
  reg [31:0] _T_4509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8624;
  reg [31:0] _T_4509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8625;
  reg [31:0] _T_4510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8626;
  reg [31:0] _T_4510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8627;
  reg [31:0] _T_4511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8628;
  reg [31:0] _T_4511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8629;
  reg [31:0] _T_4512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8630;
  reg [31:0] _T_4512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8631;
  reg [31:0] _T_4513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8632;
  reg [31:0] _T_4513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8633;
  reg [31:0] _T_4514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8634;
  reg [31:0] _T_4514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8635;
  reg [31:0] _T_4515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8636;
  reg [31:0] _T_4515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8637;
  reg [31:0] _T_4516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8638;
  reg [31:0] _T_4516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8639;
  reg [31:0] _T_4517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8640;
  reg [31:0] _T_4517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8641;
  reg [31:0] _T_4518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8642;
  reg [31:0] _T_4518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8643;
  reg [31:0] _T_4519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8644;
  reg [31:0] _T_4519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8645;
  reg [31:0] _T_4520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8646;
  reg [31:0] _T_4520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8647;
  reg [31:0] _T_4521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8648;
  reg [31:0] _T_4521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8649;
  reg [31:0] _T_4522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8650;
  reg [31:0] _T_4522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8651;
  reg [31:0] _T_4523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8652;
  reg [31:0] _T_4523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8653;
  reg [31:0] _T_4524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8654;
  reg [31:0] _T_4524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8655;
  reg [31:0] _T_4525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8656;
  reg [31:0] _T_4525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8657;
  reg [31:0] _T_4526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8658;
  reg [31:0] _T_4526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8659;
  reg [31:0] _T_4527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8660;
  reg [31:0] _T_4527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8661;
  reg [31:0] _T_4528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8662;
  reg [31:0] _T_4528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8663;
  reg [31:0] _T_4529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8664;
  reg [31:0] _T_4529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8665;
  reg [31:0] _T_4530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8666;
  reg [31:0] _T_4530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8667;
  reg [31:0] _T_4531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8668;
  reg [31:0] _T_4531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8669;
  reg [31:0] _T_4532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8670;
  reg [31:0] _T_4532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8671;
  reg [31:0] _T_4533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8672;
  reg [31:0] _T_4533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8673;
  reg [31:0] _T_4534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8674;
  reg [31:0] _T_4534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8675;
  reg [31:0] _T_4535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8676;
  reg [31:0] _T_4535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8677;
  reg [31:0] _T_4536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8678;
  reg [31:0] _T_4536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8679;
  reg [31:0] _T_4537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8680;
  reg [31:0] _T_4537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8681;
  reg [31:0] _T_4538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8682;
  reg [31:0] _T_4538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8683;
  reg [31:0] _T_4539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8684;
  reg [31:0] _T_4539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8685;
  reg [31:0] _T_4540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8686;
  reg [31:0] _T_4540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8687;
  reg [31:0] _T_4541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8688;
  reg [31:0] _T_4541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8689;
  reg [31:0] _T_4542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8690;
  reg [31:0] _T_4542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8691;
  reg [31:0] _T_4543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8692;
  reg [31:0] _T_4543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8693;
  reg [31:0] _T_4544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8694;
  reg [31:0] _T_4544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8695;
  reg [31:0] _T_4545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8696;
  reg [31:0] _T_4545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8697;
  reg [31:0] _T_4546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8698;
  reg [31:0] _T_4546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8699;
  reg [31:0] _T_4547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8700;
  reg [31:0] _T_4547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8701;
  reg [31:0] _T_4548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8702;
  reg [31:0] _T_4548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8703;
  reg [31:0] _T_4549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8704;
  reg [31:0] _T_4549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8705;
  reg [31:0] _T_4550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8706;
  reg [31:0] _T_4550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8707;
  reg [31:0] _T_4551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8708;
  reg [31:0] _T_4551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8709;
  reg [31:0] _T_4552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8710;
  reg [31:0] _T_4552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8711;
  reg [31:0] _T_4553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8712;
  reg [31:0] _T_4553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8713;
  reg [31:0] _T_4554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8714;
  reg [31:0] _T_4554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8715;
  reg [31:0] _T_4555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8716;
  reg [31:0] _T_4555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8717;
  reg [31:0] _T_4556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8718;
  reg [31:0] _T_4556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8719;
  reg [31:0] _T_4557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8720;
  reg [31:0] _T_4557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8721;
  reg [31:0] _T_4558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8722;
  reg [31:0] _T_4558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8723;
  reg [31:0] _T_4559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8724;
  reg [31:0] _T_4559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8725;
  reg [31:0] _T_4560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8726;
  reg [31:0] _T_4560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8727;
  reg [31:0] _T_4561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8728;
  reg [31:0] _T_4561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8729;
  reg [31:0] _T_4562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8730;
  reg [31:0] _T_4562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8731;
  reg [31:0] _T_4563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8732;
  reg [31:0] _T_4563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8733;
  reg [31:0] _T_4564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8734;
  reg [31:0] _T_4564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8735;
  reg [31:0] _T_4565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8736;
  reg [31:0] _T_4565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8737;
  reg [31:0] _T_4566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8738;
  reg [31:0] _T_4566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8739;
  reg [31:0] _T_4567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8740;
  reg [31:0] _T_4567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8741;
  reg [31:0] _T_4568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8742;
  reg [31:0] _T_4568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8743;
  reg [31:0] _T_4569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8744;
  reg [31:0] _T_4569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8745;
  reg [31:0] _T_4570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8746;
  reg [31:0] _T_4570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8747;
  reg [31:0] _T_4571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8748;
  reg [31:0] _T_4571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8749;
  reg [31:0] _T_4572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8750;
  reg [31:0] _T_4572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8751;
  reg [31:0] _T_4573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8752;
  reg [31:0] _T_4573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8753;
  reg [31:0] _T_4574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8754;
  reg [31:0] _T_4574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8755;
  reg [31:0] _T_4575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8756;
  reg [31:0] _T_4575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8757;
  reg [31:0] _T_4576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8758;
  reg [31:0] _T_4576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8759;
  reg [31:0] _T_4577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8760;
  reg [31:0] _T_4577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8761;
  reg [31:0] _T_4578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8762;
  reg [31:0] _T_4578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8763;
  reg [31:0] _T_4579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8764;
  reg [31:0] _T_4579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8765;
  reg [31:0] _T_4580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8766;
  reg [31:0] _T_4580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8767;
  reg [31:0] _T_4581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8768;
  reg [31:0] _T_4581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8769;
  reg [31:0] _T_4582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8770;
  reg [31:0] _T_4582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8771;
  reg [31:0] _T_4583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8772;
  reg [31:0] _T_4583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8773;
  reg [31:0] _T_4584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8774;
  reg [31:0] _T_4584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8775;
  reg [31:0] _T_4585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8776;
  reg [31:0] _T_4585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8777;
  reg [31:0] _T_4586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8778;
  reg [31:0] _T_4586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8779;
  reg [31:0] _T_4587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8780;
  reg [31:0] _T_4587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8781;
  reg [31:0] _T_4588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8782;
  reg [31:0] _T_4588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8783;
  reg [31:0] _T_4589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8784;
  reg [31:0] _T_4589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8785;
  reg [31:0] _T_4590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8786;
  reg [31:0] _T_4590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8787;
  reg [31:0] _T_4591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8788;
  reg [31:0] _T_4591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8789;
  reg [31:0] _T_4592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8790;
  reg [31:0] _T_4592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8791;
  reg [31:0] _T_4593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8792;
  reg [31:0] _T_4593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8793;
  reg [31:0] _T_4594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8794;
  reg [31:0] _T_4594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8795;
  reg [31:0] _T_4595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8796;
  reg [31:0] _T_4595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8797;
  reg [31:0] _T_4596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8798;
  reg [31:0] _T_4596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8799;
  reg [31:0] _T_4597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8800;
  reg [31:0] _T_4597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8801;
  reg [31:0] _T_4598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8802;
  reg [31:0] _T_4598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8803;
  reg [31:0] _T_4599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8804;
  reg [31:0] _T_4599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8805;
  reg [31:0] _T_4600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8806;
  reg [31:0] _T_4600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8807;
  reg [31:0] _T_4601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8808;
  reg [31:0] _T_4601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8809;
  reg [31:0] _T_4602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8810;
  reg [31:0] _T_4602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8811;
  reg [31:0] _T_4603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8812;
  reg [31:0] _T_4603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8813;
  reg [31:0] _T_4604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8814;
  reg [31:0] _T_4604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8815;
  reg [31:0] _T_4605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8816;
  reg [31:0] _T_4605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8817;
  reg [31:0] _T_4606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8818;
  reg [31:0] _T_4606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8819;
  reg [31:0] _T_4607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8820;
  reg [31:0] _T_4607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8821;
  reg [31:0] _T_4608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8822;
  reg [31:0] _T_4608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8823;
  reg [31:0] _T_4609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8824;
  reg [31:0] _T_4609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8825;
  reg [31:0] _T_4610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8826;
  reg [31:0] _T_4610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8827;
  reg [31:0] _T_4611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8828;
  reg [31:0] _T_4611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8829;
  reg [31:0] _T_4612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8830;
  reg [31:0] _T_4612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8831;
  reg [31:0] _T_4613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8832;
  reg [31:0] _T_4613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8833;
  reg [31:0] _T_4614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8834;
  reg [31:0] _T_4614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8835;
  reg [31:0] _T_4615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8836;
  reg [31:0] _T_4615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8837;
  reg [31:0] _T_4616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8838;
  reg [31:0] _T_4616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8839;
  reg [31:0] _T_4617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8840;
  reg [31:0] _T_4617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8841;
  reg [31:0] _T_4618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8842;
  reg [31:0] _T_4618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8843;
  reg [31:0] _T_4619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8844;
  reg [31:0] _T_4619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8845;
  reg [31:0] _T_4620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8846;
  reg [31:0] _T_4620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8847;
  reg [31:0] _T_4621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8848;
  reg [31:0] _T_4621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8849;
  reg [31:0] _T_4622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8850;
  reg [31:0] _T_4622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8851;
  reg [31:0] _T_4623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8852;
  reg [31:0] _T_4623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8853;
  reg [31:0] _T_4624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8854;
  reg [31:0] _T_4624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8855;
  reg [31:0] _T_4625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8856;
  reg [31:0] _T_4625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8857;
  reg [31:0] _T_4626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8858;
  reg [31:0] _T_4626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8859;
  reg [31:0] _T_4627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8860;
  reg [31:0] _T_4627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8861;
  reg [31:0] _T_4628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8862;
  reg [31:0] _T_4628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8863;
  reg [31:0] _T_4629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8864;
  reg [31:0] _T_4629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8865;
  reg [31:0] _T_4630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8866;
  reg [31:0] _T_4630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8867;
  reg [31:0] _T_4631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8868;
  reg [31:0] _T_4631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8869;
  reg [31:0] _T_4632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8870;
  reg [31:0] _T_4632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8871;
  reg [31:0] _T_4633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8872;
  reg [31:0] _T_4633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8873;
  reg [31:0] _T_4634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8874;
  reg [31:0] _T_4634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8875;
  reg [31:0] _T_4635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8876;
  reg [31:0] _T_4635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8877;
  reg [31:0] _T_4636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8878;
  reg [31:0] _T_4636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8879;
  reg [31:0] _T_4637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8880;
  reg [31:0] _T_4637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8881;
  reg [31:0] _T_4638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8882;
  reg [31:0] _T_4638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8883;
  reg [31:0] _T_4639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8884;
  reg [31:0] _T_4639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8885;
  reg [31:0] _T_4640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8886;
  reg [31:0] _T_4640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8887;
  reg [31:0] _T_4641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8888;
  reg [31:0] _T_4641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8889;
  reg [31:0] _T_4642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8890;
  reg [31:0] _T_4642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8891;
  reg [31:0] _T_4643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8892;
  reg [31:0] _T_4643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8893;
  reg [31:0] _T_4644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8894;
  reg [31:0] _T_4644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8895;
  reg [31:0] _T_4645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8896;
  reg [31:0] _T_4645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8897;
  reg [31:0] _T_4646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8898;
  reg [31:0] _T_4646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8899;
  reg [31:0] _T_4647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8900;
  reg [31:0] _T_4647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8901;
  reg [31:0] _T_4648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8902;
  reg [31:0] _T_4648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8903;
  reg [31:0] _T_4649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8904;
  reg [31:0] _T_4649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8905;
  reg [31:0] _T_4650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8906;
  reg [31:0] _T_4650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8907;
  reg [31:0] _T_4651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8908;
  reg [31:0] _T_4651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8909;
  reg [31:0] _T_4652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8910;
  reg [31:0] _T_4652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8911;
  reg [31:0] _T_4653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8912;
  reg [31:0] _T_4653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8913;
  reg [31:0] _T_4654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8914;
  reg [31:0] _T_4654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8915;
  reg [31:0] _T_4655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8916;
  reg [31:0] _T_4655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8917;
  reg [31:0] _T_4656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8918;
  reg [31:0] _T_4656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8919;
  reg [31:0] _T_4657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8920;
  reg [31:0] _T_4657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8921;
  reg [31:0] _T_4658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8922;
  reg [31:0] _T_4658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8923;
  reg [31:0] _T_4659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8924;
  reg [31:0] _T_4659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8925;
  reg [31:0] _T_4660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8926;
  reg [31:0] _T_4660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8927;
  reg [31:0] _T_4661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8928;
  reg [31:0] _T_4661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8929;
  reg [31:0] _T_4662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8930;
  reg [31:0] _T_4662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8931;
  reg [31:0] _T_4663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8932;
  reg [31:0] _T_4663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8933;
  reg [31:0] _T_4664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8934;
  reg [31:0] _T_4664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8935;
  reg [31:0] _T_4665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8936;
  reg [31:0] _T_4665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8937;
  reg [31:0] _T_4666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8938;
  reg [31:0] _T_4666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8939;
  reg [31:0] _T_4667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8940;
  reg [31:0] _T_4667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8941;
  reg [31:0] _T_4668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8942;
  reg [31:0] _T_4668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8943;
  reg [31:0] _T_4669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8944;
  reg [31:0] _T_4669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8945;
  reg [31:0] _T_4670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8946;
  reg [31:0] _T_4670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8947;
  reg [31:0] _T_4671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8948;
  reg [31:0] _T_4671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8949;
  reg [31:0] _T_4672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8950;
  reg [31:0] _T_4672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8951;
  reg [31:0] _T_4673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8952;
  reg [31:0] _T_4673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8953;
  reg [31:0] _T_4674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8954;
  reg [31:0] _T_4674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8955;
  reg [31:0] _T_4675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8956;
  reg [31:0] _T_4675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8957;
  reg [31:0] _T_4676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8958;
  reg [31:0] _T_4676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8959;
  reg [31:0] _T_4677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8960;
  reg [31:0] _T_4677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8961;
  reg [31:0] _T_4678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8962;
  reg [31:0] _T_4678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8963;
  reg [31:0] _T_4679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8964;
  reg [31:0] _T_4679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8965;
  reg [31:0] _T_4680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8966;
  reg [31:0] _T_4680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8967;
  reg [31:0] _T_4681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8968;
  reg [31:0] _T_4681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8969;
  reg [31:0] _T_4682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8970;
  reg [31:0] _T_4682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8971;
  reg [31:0] _T_4683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8972;
  reg [31:0] _T_4683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8973;
  reg [31:0] _T_4684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8974;
  reg [31:0] _T_4684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8975;
  reg [31:0] _T_4685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8976;
  reg [31:0] _T_4685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8977;
  reg [31:0] _T_4686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8978;
  reg [31:0] _T_4686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8979;
  reg [31:0] _T_4687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8980;
  reg [31:0] _T_4687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8981;
  reg [31:0] _T_4688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8982;
  reg [31:0] _T_4688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8983;
  reg [31:0] _T_4689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8984;
  reg [31:0] _T_4689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8985;
  reg [31:0] _T_4690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8986;
  reg [31:0] _T_4690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8987;
  reg [31:0] _T_4691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8988;
  reg [31:0] _T_4691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8989;
  reg [31:0] _T_4692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8990;
  reg [31:0] _T_4692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8991;
  reg [31:0] _T_4693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8992;
  reg [31:0] _T_4693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8993;
  reg [31:0] _T_4694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8994;
  reg [31:0] _T_4694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8995;
  reg [31:0] _T_4695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8996;
  reg [31:0] _T_4695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8997;
  reg [31:0] _T_4696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8998;
  reg [31:0] _T_4696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8999;
  reg [31:0] _T_4697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9000;
  reg [31:0] _T_4697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9001;
  reg [31:0] _T_4698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9002;
  reg [31:0] _T_4698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9003;
  reg [31:0] _T_4699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9004;
  reg [31:0] _T_4699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9005;
  reg [31:0] _T_4700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9006;
  reg [31:0] _T_4700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9007;
  reg [31:0] _T_4701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9008;
  reg [31:0] _T_4701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9009;
  reg [31:0] _T_4702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9010;
  reg [31:0] _T_4702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9011;
  reg [31:0] _T_4703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9012;
  reg [31:0] _T_4703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9013;
  reg [31:0] _T_4704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9014;
  reg [31:0] _T_4704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9015;
  reg [31:0] _T_4705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9016;
  reg [31:0] _T_4705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9017;
  reg [31:0] _T_4706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9018;
  reg [31:0] _T_4706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9019;
  reg [31:0] _T_4707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9020;
  reg [31:0] _T_4707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9021;
  reg [31:0] _T_4708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9022;
  reg [31:0] _T_4708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9023;
  reg [31:0] _T_4709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9024;
  reg [31:0] _T_4709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9025;
  reg [31:0] _T_4710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9026;
  reg [31:0] _T_4710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9027;
  reg [31:0] _T_4711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9028;
  reg [31:0] _T_4711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9029;
  reg [31:0] _T_4712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9030;
  reg [31:0] _T_4712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9031;
  reg [31:0] _T_4713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9032;
  reg [31:0] _T_4713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9033;
  reg [31:0] _T_4714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9034;
  reg [31:0] _T_4714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9035;
  reg [31:0] _T_4715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9036;
  reg [31:0] _T_4715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9037;
  reg [31:0] _T_4716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9038;
  reg [31:0] _T_4716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9039;
  reg [31:0] _T_4717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9040;
  reg [31:0] _T_4717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9041;
  reg [31:0] _T_4718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9042;
  reg [31:0] _T_4718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9043;
  reg [31:0] _T_4719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9044;
  reg [31:0] _T_4719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9045;
  reg [31:0] _T_4720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9046;
  reg [31:0] _T_4720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9047;
  reg [31:0] _T_4721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9048;
  reg [31:0] _T_4721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9049;
  reg [31:0] _T_4722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9050;
  reg [31:0] _T_4722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9051;
  reg [31:0] _T_4723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9052;
  reg [31:0] _T_4723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9053;
  reg [31:0] _T_4724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9054;
  reg [31:0] _T_4724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9055;
  reg [31:0] _T_4725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9056;
  reg [31:0] _T_4725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9057;
  reg [31:0] _T_4726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9058;
  reg [31:0] _T_4726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9059;
  reg [31:0] _T_4727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9060;
  reg [31:0] _T_4727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9061;
  reg [31:0] _T_4728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9062;
  reg [31:0] _T_4728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9063;
  reg [31:0] _T_4729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9064;
  reg [31:0] _T_4729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9065;
  reg [31:0] _T_4730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9066;
  reg [31:0] _T_4730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9067;
  reg [31:0] _T_4731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9068;
  reg [31:0] _T_4731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9069;
  reg [31:0] _T_4732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9070;
  reg [31:0] _T_4732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9071;
  reg [31:0] _T_4733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9072;
  reg [31:0] _T_4733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9073;
  reg [31:0] _T_4734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9074;
  reg [31:0] _T_4734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9075;
  reg [31:0] _T_4735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9076;
  reg [31:0] _T_4735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9077;
  reg [31:0] _T_4736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9078;
  reg [31:0] _T_4736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9079;
  reg [31:0] _T_4737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9080;
  reg [31:0] _T_4737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9081;
  reg [31:0] _T_4738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9082;
  reg [31:0] _T_4738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9083;
  reg [31:0] _T_4739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9084;
  reg [31:0] _T_4739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9085;
  reg [31:0] _T_4740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9086;
  reg [31:0] _T_4740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9087;
  reg [31:0] _T_4741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9088;
  reg [31:0] _T_4741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9089;
  reg [31:0] _T_4742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9090;
  reg [31:0] _T_4742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9091;
  reg [31:0] _T_4743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9092;
  reg [31:0] _T_4743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9093;
  reg [31:0] _T_4744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9094;
  reg [31:0] _T_4744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9095;
  reg [31:0] _T_4745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9096;
  reg [31:0] _T_4745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9097;
  reg [31:0] _T_4746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9098;
  reg [31:0] _T_4746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9099;
  reg [31:0] _T_4747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9100;
  reg [31:0] _T_4747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9101;
  reg [31:0] _T_4748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9102;
  reg [31:0] _T_4748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9103;
  reg [31:0] _T_4749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9104;
  reg [31:0] _T_4749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9105;
  reg [31:0] _T_4750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9106;
  reg [31:0] _T_4750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9107;
  reg [31:0] _T_4751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9108;
  reg [31:0] _T_4751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9109;
  reg [31:0] _T_4752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9110;
  reg [31:0] _T_4752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9111;
  reg [31:0] _T_4753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9112;
  reg [31:0] _T_4753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9113;
  reg [31:0] _T_4754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9114;
  reg [31:0] _T_4754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9115;
  reg [31:0] _T_4755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9116;
  reg [31:0] _T_4755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9117;
  reg [31:0] _T_4756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9118;
  reg [31:0] _T_4756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9119;
  reg [31:0] _T_4757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9120;
  reg [31:0] _T_4757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9121;
  reg [31:0] _T_4758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9122;
  reg [31:0] _T_4758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9123;
  reg [31:0] _T_4759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9124;
  reg [31:0] _T_4759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9125;
  reg [31:0] _T_4760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9126;
  reg [31:0] _T_4760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9127;
  reg [31:0] _T_4761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9128;
  reg [31:0] _T_4761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9129;
  reg [31:0] _T_4762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9130;
  reg [31:0] _T_4762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9131;
  reg [31:0] _T_4763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9132;
  reg [31:0] _T_4763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9133;
  reg [31:0] _T_4764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9134;
  reg [31:0] _T_4764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9135;
  reg [31:0] _T_4765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9136;
  reg [31:0] _T_4765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9137;
  reg [31:0] _T_4766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9138;
  reg [31:0] _T_4766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9139;
  reg [31:0] _T_4767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9140;
  reg [31:0] _T_4767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9141;
  reg [31:0] _T_4768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9142;
  reg [31:0] _T_4768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9143;
  reg [31:0] _T_4769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9144;
  reg [31:0] _T_4769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9145;
  reg [31:0] _T_4770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9146;
  reg [31:0] _T_4770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9147;
  reg [31:0] _T_4771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9148;
  reg [31:0] _T_4771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9149;
  reg [31:0] _T_4772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9150;
  reg [31:0] _T_4772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9151;
  reg [31:0] _T_4773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9152;
  reg [31:0] _T_4773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9153;
  reg [31:0] _T_4774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9154;
  reg [31:0] _T_4774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9155;
  reg [31:0] _T_4775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9156;
  reg [31:0] _T_4775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9157;
  reg [31:0] _T_4776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9158;
  reg [31:0] _T_4776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9159;
  reg [31:0] _T_4777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9160;
  reg [31:0] _T_4777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9161;
  reg [31:0] _T_4778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9162;
  reg [31:0] _T_4778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9163;
  reg [31:0] _T_4779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9164;
  reg [31:0] _T_4779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9165;
  reg [31:0] _T_4780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9166;
  reg [31:0] _T_4780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9167;
  reg [31:0] _T_4781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9168;
  reg [31:0] _T_4781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9169;
  reg [31:0] _T_4782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9170;
  reg [31:0] _T_4782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9171;
  reg [31:0] _T_4783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9172;
  reg [31:0] _T_4783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9173;
  reg [31:0] _T_4784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9174;
  reg [31:0] _T_4784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9175;
  reg [31:0] _T_4785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9176;
  reg [31:0] _T_4785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9177;
  reg [31:0] _T_4786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9178;
  reg [31:0] _T_4786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9179;
  reg [31:0] _T_4787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9180;
  reg [31:0] _T_4787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9181;
  reg [31:0] _T_4788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9182;
  reg [31:0] _T_4788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9183;
  reg [31:0] _T_4789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9184;
  reg [31:0] _T_4789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9185;
  reg [31:0] _T_4790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9186;
  reg [31:0] _T_4790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9187;
  reg [31:0] _T_4791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9188;
  reg [31:0] _T_4791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9189;
  reg [31:0] _T_4792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9190;
  reg [31:0] _T_4792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9191;
  reg [31:0] _T_4793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9192;
  reg [31:0] _T_4793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9193;
  reg [31:0] _T_4794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9194;
  reg [31:0] _T_4794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9195;
  reg [31:0] _T_4795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9196;
  reg [31:0] _T_4795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9197;
  reg [31:0] _T_4796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9198;
  reg [31:0] _T_4796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9199;
  reg [31:0] _T_4797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9200;
  reg [31:0] _T_4797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9201;
  reg [31:0] _T_4798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9202;
  reg [31:0] _T_4798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9203;
  reg [31:0] _T_4799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9204;
  reg [31:0] _T_4799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9205;
  reg [31:0] _T_4800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9206;
  reg [31:0] _T_4800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9207;
  reg [31:0] _T_4801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9208;
  reg [31:0] _T_4801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9209;
  reg [31:0] _T_4802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9210;
  reg [31:0] _T_4802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9211;
  reg [31:0] _T_4803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9212;
  reg [31:0] _T_4803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9213;
  reg [31:0] _T_4804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9214;
  reg [31:0] _T_4804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9215;
  reg [31:0] _T_4805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9216;
  reg [31:0] _T_4805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9217;
  wire [31:0] _GEN_15362 = 9'h1 == cnt[8:0] ? $signed(32'shffff) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15363 = 9'h2 == cnt[8:0] ? $signed(32'shfffb) : $signed(_GEN_15362); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15364 = 9'h3 == cnt[8:0] ? $signed(32'shfff5) : $signed(_GEN_15363); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15365 = 9'h4 == cnt[8:0] ? $signed(32'shffec) : $signed(_GEN_15364); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15366 = 9'h5 == cnt[8:0] ? $signed(32'shffe1) : $signed(_GEN_15365); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15367 = 9'h6 == cnt[8:0] ? $signed(32'shffd4) : $signed(_GEN_15366); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15368 = 9'h7 == cnt[8:0] ? $signed(32'shffc4) : $signed(_GEN_15367); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15369 = 9'h8 == cnt[8:0] ? $signed(32'shffb1) : $signed(_GEN_15368); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15370 = 9'h9 == cnt[8:0] ? $signed(32'shff9c) : $signed(_GEN_15369); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15371 = 9'ha == cnt[8:0] ? $signed(32'shff85) : $signed(_GEN_15370); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15372 = 9'hb == cnt[8:0] ? $signed(32'shff6b) : $signed(_GEN_15371); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15373 = 9'hc == cnt[8:0] ? $signed(32'shff4e) : $signed(_GEN_15372); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15374 = 9'hd == cnt[8:0] ? $signed(32'shff30) : $signed(_GEN_15373); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15375 = 9'he == cnt[8:0] ? $signed(32'shff0e) : $signed(_GEN_15374); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15376 = 9'hf == cnt[8:0] ? $signed(32'shfeeb) : $signed(_GEN_15375); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15377 = 9'h10 == cnt[8:0] ? $signed(32'shfec4) : $signed(_GEN_15376); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15378 = 9'h11 == cnt[8:0] ? $signed(32'shfe9c) : $signed(_GEN_15377); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15379 = 9'h12 == cnt[8:0] ? $signed(32'shfe71) : $signed(_GEN_15378); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15380 = 9'h13 == cnt[8:0] ? $signed(32'shfe43) : $signed(_GEN_15379); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15381 = 9'h14 == cnt[8:0] ? $signed(32'shfe13) : $signed(_GEN_15380); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15382 = 9'h15 == cnt[8:0] ? $signed(32'shfde1) : $signed(_GEN_15381); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15383 = 9'h16 == cnt[8:0] ? $signed(32'shfdac) : $signed(_GEN_15382); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15384 = 9'h17 == cnt[8:0] ? $signed(32'shfd74) : $signed(_GEN_15383); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15385 = 9'h18 == cnt[8:0] ? $signed(32'shfd3b) : $signed(_GEN_15384); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15386 = 9'h19 == cnt[8:0] ? $signed(32'shfcfe) : $signed(_GEN_15385); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15387 = 9'h1a == cnt[8:0] ? $signed(32'shfcc0) : $signed(_GEN_15386); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15388 = 9'h1b == cnt[8:0] ? $signed(32'shfc7f) : $signed(_GEN_15387); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15389 = 9'h1c == cnt[8:0] ? $signed(32'shfc3b) : $signed(_GEN_15388); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15390 = 9'h1d == cnt[8:0] ? $signed(32'shfbf5) : $signed(_GEN_15389); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15391 = 9'h1e == cnt[8:0] ? $signed(32'shfbad) : $signed(_GEN_15390); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15392 = 9'h1f == cnt[8:0] ? $signed(32'shfb62) : $signed(_GEN_15391); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15393 = 9'h20 == cnt[8:0] ? $signed(32'shfb15) : $signed(_GEN_15392); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15394 = 9'h21 == cnt[8:0] ? $signed(32'shfac5) : $signed(_GEN_15393); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15395 = 9'h22 == cnt[8:0] ? $signed(32'shfa73) : $signed(_GEN_15394); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15396 = 9'h23 == cnt[8:0] ? $signed(32'shfa1f) : $signed(_GEN_15395); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15397 = 9'h24 == cnt[8:0] ? $signed(32'shf9c8) : $signed(_GEN_15396); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15398 = 9'h25 == cnt[8:0] ? $signed(32'shf96e) : $signed(_GEN_15397); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15399 = 9'h26 == cnt[8:0] ? $signed(32'shf913) : $signed(_GEN_15398); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15400 = 9'h27 == cnt[8:0] ? $signed(32'shf8b4) : $signed(_GEN_15399); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15401 = 9'h28 == cnt[8:0] ? $signed(32'shf854) : $signed(_GEN_15400); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15402 = 9'h29 == cnt[8:0] ? $signed(32'shf7f1) : $signed(_GEN_15401); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15403 = 9'h2a == cnt[8:0] ? $signed(32'shf78c) : $signed(_GEN_15402); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15404 = 9'h2b == cnt[8:0] ? $signed(32'shf724) : $signed(_GEN_15403); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15405 = 9'h2c == cnt[8:0] ? $signed(32'shf6ba) : $signed(_GEN_15404); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15406 = 9'h2d == cnt[8:0] ? $signed(32'shf64e) : $signed(_GEN_15405); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15407 = 9'h2e == cnt[8:0] ? $signed(32'shf5df) : $signed(_GEN_15406); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15408 = 9'h2f == cnt[8:0] ? $signed(32'shf56e) : $signed(_GEN_15407); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15409 = 9'h30 == cnt[8:0] ? $signed(32'shf4fa) : $signed(_GEN_15408); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15410 = 9'h31 == cnt[8:0] ? $signed(32'shf484) : $signed(_GEN_15409); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15411 = 9'h32 == cnt[8:0] ? $signed(32'shf40c) : $signed(_GEN_15410); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15412 = 9'h33 == cnt[8:0] ? $signed(32'shf391) : $signed(_GEN_15411); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15413 = 9'h34 == cnt[8:0] ? $signed(32'shf314) : $signed(_GEN_15412); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15414 = 9'h35 == cnt[8:0] ? $signed(32'shf295) : $signed(_GEN_15413); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15415 = 9'h36 == cnt[8:0] ? $signed(32'shf213) : $signed(_GEN_15414); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15416 = 9'h37 == cnt[8:0] ? $signed(32'shf18f) : $signed(_GEN_15415); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15417 = 9'h38 == cnt[8:0] ? $signed(32'shf109) : $signed(_GEN_15416); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15418 = 9'h39 == cnt[8:0] ? $signed(32'shf080) : $signed(_GEN_15417); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15419 = 9'h3a == cnt[8:0] ? $signed(32'sheff5) : $signed(_GEN_15418); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15420 = 9'h3b == cnt[8:0] ? $signed(32'shef68) : $signed(_GEN_15419); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15421 = 9'h3c == cnt[8:0] ? $signed(32'sheed9) : $signed(_GEN_15420); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15422 = 9'h3d == cnt[8:0] ? $signed(32'shee47) : $signed(_GEN_15421); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15423 = 9'h3e == cnt[8:0] ? $signed(32'shedb3) : $signed(_GEN_15422); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15424 = 9'h3f == cnt[8:0] ? $signed(32'shed1c) : $signed(_GEN_15423); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15425 = 9'h40 == cnt[8:0] ? $signed(32'shec83) : $signed(_GEN_15424); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15426 = 9'h41 == cnt[8:0] ? $signed(32'shebe8) : $signed(_GEN_15425); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15427 = 9'h42 == cnt[8:0] ? $signed(32'sheb4b) : $signed(_GEN_15426); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15428 = 9'h43 == cnt[8:0] ? $signed(32'sheaab) : $signed(_GEN_15427); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15429 = 9'h44 == cnt[8:0] ? $signed(32'shea0a) : $signed(_GEN_15428); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15430 = 9'h45 == cnt[8:0] ? $signed(32'she966) : $signed(_GEN_15429); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15431 = 9'h46 == cnt[8:0] ? $signed(32'she8bf) : $signed(_GEN_15430); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15432 = 9'h47 == cnt[8:0] ? $signed(32'she817) : $signed(_GEN_15431); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15433 = 9'h48 == cnt[8:0] ? $signed(32'she76c) : $signed(_GEN_15432); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15434 = 9'h49 == cnt[8:0] ? $signed(32'she6bf) : $signed(_GEN_15433); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15435 = 9'h4a == cnt[8:0] ? $signed(32'she610) : $signed(_GEN_15434); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15436 = 9'h4b == cnt[8:0] ? $signed(32'she55e) : $signed(_GEN_15435); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15437 = 9'h4c == cnt[8:0] ? $signed(32'she4aa) : $signed(_GEN_15436); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15438 = 9'h4d == cnt[8:0] ? $signed(32'she3f4) : $signed(_GEN_15437); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15439 = 9'h4e == cnt[8:0] ? $signed(32'she33c) : $signed(_GEN_15438); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15440 = 9'h4f == cnt[8:0] ? $signed(32'she282) : $signed(_GEN_15439); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15441 = 9'h50 == cnt[8:0] ? $signed(32'she1c6) : $signed(_GEN_15440); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15442 = 9'h51 == cnt[8:0] ? $signed(32'she107) : $signed(_GEN_15441); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15443 = 9'h52 == cnt[8:0] ? $signed(32'she046) : $signed(_GEN_15442); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15444 = 9'h53 == cnt[8:0] ? $signed(32'shdf83) : $signed(_GEN_15443); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15445 = 9'h54 == cnt[8:0] ? $signed(32'shdebe) : $signed(_GEN_15444); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15446 = 9'h55 == cnt[8:0] ? $signed(32'shddf7) : $signed(_GEN_15445); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15447 = 9'h56 == cnt[8:0] ? $signed(32'shdd2d) : $signed(_GEN_15446); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15448 = 9'h57 == cnt[8:0] ? $signed(32'shdc62) : $signed(_GEN_15447); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15449 = 9'h58 == cnt[8:0] ? $signed(32'shdb94) : $signed(_GEN_15448); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15450 = 9'h59 == cnt[8:0] ? $signed(32'shdac4) : $signed(_GEN_15449); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15451 = 9'h5a == cnt[8:0] ? $signed(32'shd9f2) : $signed(_GEN_15450); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15452 = 9'h5b == cnt[8:0] ? $signed(32'shd91e) : $signed(_GEN_15451); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15453 = 9'h5c == cnt[8:0] ? $signed(32'shd848) : $signed(_GEN_15452); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15454 = 9'h5d == cnt[8:0] ? $signed(32'shd770) : $signed(_GEN_15453); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15455 = 9'h5e == cnt[8:0] ? $signed(32'shd696) : $signed(_GEN_15454); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15456 = 9'h5f == cnt[8:0] ? $signed(32'shd5ba) : $signed(_GEN_15455); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15457 = 9'h60 == cnt[8:0] ? $signed(32'shd4db) : $signed(_GEN_15456); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15458 = 9'h61 == cnt[8:0] ? $signed(32'shd3fb) : $signed(_GEN_15457); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15459 = 9'h62 == cnt[8:0] ? $signed(32'shd318) : $signed(_GEN_15458); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15460 = 9'h63 == cnt[8:0] ? $signed(32'shd234) : $signed(_GEN_15459); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15461 = 9'h64 == cnt[8:0] ? $signed(32'shd14d) : $signed(_GEN_15460); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15462 = 9'h65 == cnt[8:0] ? $signed(32'shd065) : $signed(_GEN_15461); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15463 = 9'h66 == cnt[8:0] ? $signed(32'shcf7a) : $signed(_GEN_15462); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15464 = 9'h67 == cnt[8:0] ? $signed(32'shce8e) : $signed(_GEN_15463); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15465 = 9'h68 == cnt[8:0] ? $signed(32'shcd9f) : $signed(_GEN_15464); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15466 = 9'h69 == cnt[8:0] ? $signed(32'shccae) : $signed(_GEN_15465); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15467 = 9'h6a == cnt[8:0] ? $signed(32'shcbbc) : $signed(_GEN_15466); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15468 = 9'h6b == cnt[8:0] ? $signed(32'shcac7) : $signed(_GEN_15467); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15469 = 9'h6c == cnt[8:0] ? $signed(32'shc9d1) : $signed(_GEN_15468); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15470 = 9'h6d == cnt[8:0] ? $signed(32'shc8d9) : $signed(_GEN_15469); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15471 = 9'h6e == cnt[8:0] ? $signed(32'shc7de) : $signed(_GEN_15470); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15472 = 9'h6f == cnt[8:0] ? $signed(32'shc6e2) : $signed(_GEN_15471); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15473 = 9'h70 == cnt[8:0] ? $signed(32'shc5e4) : $signed(_GEN_15472); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15474 = 9'h71 == cnt[8:0] ? $signed(32'shc4e4) : $signed(_GEN_15473); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15475 = 9'h72 == cnt[8:0] ? $signed(32'shc3e2) : $signed(_GEN_15474); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15476 = 9'h73 == cnt[8:0] ? $signed(32'shc2de) : $signed(_GEN_15475); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15477 = 9'h74 == cnt[8:0] ? $signed(32'shc1d8) : $signed(_GEN_15476); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15478 = 9'h75 == cnt[8:0] ? $signed(32'shc0d1) : $signed(_GEN_15477); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15479 = 9'h76 == cnt[8:0] ? $signed(32'shbfc7) : $signed(_GEN_15478); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15480 = 9'h77 == cnt[8:0] ? $signed(32'shbebc) : $signed(_GEN_15479); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15481 = 9'h78 == cnt[8:0] ? $signed(32'shbdaf) : $signed(_GEN_15480); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15482 = 9'h79 == cnt[8:0] ? $signed(32'shbca0) : $signed(_GEN_15481); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15483 = 9'h7a == cnt[8:0] ? $signed(32'shbb8f) : $signed(_GEN_15482); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15484 = 9'h7b == cnt[8:0] ? $signed(32'shba7d) : $signed(_GEN_15483); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15485 = 9'h7c == cnt[8:0] ? $signed(32'shb968) : $signed(_GEN_15484); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15486 = 9'h7d == cnt[8:0] ? $signed(32'shb852) : $signed(_GEN_15485); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15487 = 9'h7e == cnt[8:0] ? $signed(32'shb73a) : $signed(_GEN_15486); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15488 = 9'h7f == cnt[8:0] ? $signed(32'shb620) : $signed(_GEN_15487); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15489 = 9'h80 == cnt[8:0] ? $signed(32'shb505) : $signed(_GEN_15488); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15490 = 9'h81 == cnt[8:0] ? $signed(32'shb3e8) : $signed(_GEN_15489); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15491 = 9'h82 == cnt[8:0] ? $signed(32'shb2c9) : $signed(_GEN_15490); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15492 = 9'h83 == cnt[8:0] ? $signed(32'shb1a8) : $signed(_GEN_15491); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15493 = 9'h84 == cnt[8:0] ? $signed(32'shb086) : $signed(_GEN_15492); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15494 = 9'h85 == cnt[8:0] ? $signed(32'shaf62) : $signed(_GEN_15493); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15495 = 9'h86 == cnt[8:0] ? $signed(32'shae3c) : $signed(_GEN_15494); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15496 = 9'h87 == cnt[8:0] ? $signed(32'shad14) : $signed(_GEN_15495); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15497 = 9'h88 == cnt[8:0] ? $signed(32'shabeb) : $signed(_GEN_15496); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15498 = 9'h89 == cnt[8:0] ? $signed(32'shaac1) : $signed(_GEN_15497); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15499 = 9'h8a == cnt[8:0] ? $signed(32'sha994) : $signed(_GEN_15498); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15500 = 9'h8b == cnt[8:0] ? $signed(32'sha866) : $signed(_GEN_15499); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15501 = 9'h8c == cnt[8:0] ? $signed(32'sha736) : $signed(_GEN_15500); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15502 = 9'h8d == cnt[8:0] ? $signed(32'sha605) : $signed(_GEN_15501); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15503 = 9'h8e == cnt[8:0] ? $signed(32'sha4d2) : $signed(_GEN_15502); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15504 = 9'h8f == cnt[8:0] ? $signed(32'sha39e) : $signed(_GEN_15503); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15505 = 9'h90 == cnt[8:0] ? $signed(32'sha268) : $signed(_GEN_15504); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15506 = 9'h91 == cnt[8:0] ? $signed(32'sha130) : $signed(_GEN_15505); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15507 = 9'h92 == cnt[8:0] ? $signed(32'sh9ff7) : $signed(_GEN_15506); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15508 = 9'h93 == cnt[8:0] ? $signed(32'sh9ebc) : $signed(_GEN_15507); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15509 = 9'h94 == cnt[8:0] ? $signed(32'sh9d80) : $signed(_GEN_15508); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15510 = 9'h95 == cnt[8:0] ? $signed(32'sh9c42) : $signed(_GEN_15509); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15511 = 9'h96 == cnt[8:0] ? $signed(32'sh9b03) : $signed(_GEN_15510); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15512 = 9'h97 == cnt[8:0] ? $signed(32'sh99c2) : $signed(_GEN_15511); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15513 = 9'h98 == cnt[8:0] ? $signed(32'sh9880) : $signed(_GEN_15512); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15514 = 9'h99 == cnt[8:0] ? $signed(32'sh973c) : $signed(_GEN_15513); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15515 = 9'h9a == cnt[8:0] ? $signed(32'sh95f7) : $signed(_GEN_15514); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15516 = 9'h9b == cnt[8:0] ? $signed(32'sh94b0) : $signed(_GEN_15515); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15517 = 9'h9c == cnt[8:0] ? $signed(32'sh9368) : $signed(_GEN_15516); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15518 = 9'h9d == cnt[8:0] ? $signed(32'sh921f) : $signed(_GEN_15517); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15519 = 9'h9e == cnt[8:0] ? $signed(32'sh90d4) : $signed(_GEN_15518); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15520 = 9'h9f == cnt[8:0] ? $signed(32'sh8f88) : $signed(_GEN_15519); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15521 = 9'ha0 == cnt[8:0] ? $signed(32'sh8e3a) : $signed(_GEN_15520); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15522 = 9'ha1 == cnt[8:0] ? $signed(32'sh8ceb) : $signed(_GEN_15521); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15523 = 9'ha2 == cnt[8:0] ? $signed(32'sh8b9a) : $signed(_GEN_15522); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15524 = 9'ha3 == cnt[8:0] ? $signed(32'sh8a49) : $signed(_GEN_15523); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15525 = 9'ha4 == cnt[8:0] ? $signed(32'sh88f6) : $signed(_GEN_15524); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15526 = 9'ha5 == cnt[8:0] ? $signed(32'sh87a1) : $signed(_GEN_15525); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15527 = 9'ha6 == cnt[8:0] ? $signed(32'sh864c) : $signed(_GEN_15526); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15528 = 9'ha7 == cnt[8:0] ? $signed(32'sh84f5) : $signed(_GEN_15527); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15529 = 9'ha8 == cnt[8:0] ? $signed(32'sh839c) : $signed(_GEN_15528); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15530 = 9'ha9 == cnt[8:0] ? $signed(32'sh8243) : $signed(_GEN_15529); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15531 = 9'haa == cnt[8:0] ? $signed(32'sh80e8) : $signed(_GEN_15530); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15532 = 9'hab == cnt[8:0] ? $signed(32'sh7f8c) : $signed(_GEN_15531); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15533 = 9'hac == cnt[8:0] ? $signed(32'sh7e2f) : $signed(_GEN_15532); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15534 = 9'had == cnt[8:0] ? $signed(32'sh7cd0) : $signed(_GEN_15533); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15535 = 9'hae == cnt[8:0] ? $signed(32'sh7b70) : $signed(_GEN_15534); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15536 = 9'haf == cnt[8:0] ? $signed(32'sh7a10) : $signed(_GEN_15535); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15537 = 9'hb0 == cnt[8:0] ? $signed(32'sh78ad) : $signed(_GEN_15536); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15538 = 9'hb1 == cnt[8:0] ? $signed(32'sh774a) : $signed(_GEN_15537); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15539 = 9'hb2 == cnt[8:0] ? $signed(32'sh75e6) : $signed(_GEN_15538); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15540 = 9'hb3 == cnt[8:0] ? $signed(32'sh7480) : $signed(_GEN_15539); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15541 = 9'hb4 == cnt[8:0] ? $signed(32'sh731a) : $signed(_GEN_15540); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15542 = 9'hb5 == cnt[8:0] ? $signed(32'sh71b2) : $signed(_GEN_15541); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15543 = 9'hb6 == cnt[8:0] ? $signed(32'sh7049) : $signed(_GEN_15542); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15544 = 9'hb7 == cnt[8:0] ? $signed(32'sh6edf) : $signed(_GEN_15543); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15545 = 9'hb8 == cnt[8:0] ? $signed(32'sh6d74) : $signed(_GEN_15544); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15546 = 9'hb9 == cnt[8:0] ? $signed(32'sh6c08) : $signed(_GEN_15545); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15547 = 9'hba == cnt[8:0] ? $signed(32'sh6a9b) : $signed(_GEN_15546); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15548 = 9'hbb == cnt[8:0] ? $signed(32'sh692d) : $signed(_GEN_15547); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15549 = 9'hbc == cnt[8:0] ? $signed(32'sh67be) : $signed(_GEN_15548); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15550 = 9'hbd == cnt[8:0] ? $signed(32'sh664e) : $signed(_GEN_15549); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15551 = 9'hbe == cnt[8:0] ? $signed(32'sh64dd) : $signed(_GEN_15550); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15552 = 9'hbf == cnt[8:0] ? $signed(32'sh636b) : $signed(_GEN_15551); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15553 = 9'hc0 == cnt[8:0] ? $signed(32'sh61f8) : $signed(_GEN_15552); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15554 = 9'hc1 == cnt[8:0] ? $signed(32'sh6084) : $signed(_GEN_15553); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15555 = 9'hc2 == cnt[8:0] ? $signed(32'sh5f0f) : $signed(_GEN_15554); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15556 = 9'hc3 == cnt[8:0] ? $signed(32'sh5d99) : $signed(_GEN_15555); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15557 = 9'hc4 == cnt[8:0] ? $signed(32'sh5c22) : $signed(_GEN_15556); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15558 = 9'hc5 == cnt[8:0] ? $signed(32'sh5aaa) : $signed(_GEN_15557); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15559 = 9'hc6 == cnt[8:0] ? $signed(32'sh5932) : $signed(_GEN_15558); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15560 = 9'hc7 == cnt[8:0] ? $signed(32'sh57b9) : $signed(_GEN_15559); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15561 = 9'hc8 == cnt[8:0] ? $signed(32'sh563e) : $signed(_GEN_15560); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15562 = 9'hc9 == cnt[8:0] ? $signed(32'sh54c3) : $signed(_GEN_15561); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15563 = 9'hca == cnt[8:0] ? $signed(32'sh5348) : $signed(_GEN_15562); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15564 = 9'hcb == cnt[8:0] ? $signed(32'sh51cb) : $signed(_GEN_15563); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15565 = 9'hcc == cnt[8:0] ? $signed(32'sh504d) : $signed(_GEN_15564); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15566 = 9'hcd == cnt[8:0] ? $signed(32'sh4ecf) : $signed(_GEN_15565); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15567 = 9'hce == cnt[8:0] ? $signed(32'sh4d50) : $signed(_GEN_15566); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15568 = 9'hcf == cnt[8:0] ? $signed(32'sh4bd1) : $signed(_GEN_15567); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15569 = 9'hd0 == cnt[8:0] ? $signed(32'sh4a50) : $signed(_GEN_15568); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15570 = 9'hd1 == cnt[8:0] ? $signed(32'sh48cf) : $signed(_GEN_15569); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15571 = 9'hd2 == cnt[8:0] ? $signed(32'sh474d) : $signed(_GEN_15570); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15572 = 9'hd3 == cnt[8:0] ? $signed(32'sh45cb) : $signed(_GEN_15571); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15573 = 9'hd4 == cnt[8:0] ? $signed(32'sh4447) : $signed(_GEN_15572); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15574 = 9'hd5 == cnt[8:0] ? $signed(32'sh42c3) : $signed(_GEN_15573); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15575 = 9'hd6 == cnt[8:0] ? $signed(32'sh413f) : $signed(_GEN_15574); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15576 = 9'hd7 == cnt[8:0] ? $signed(32'sh3fba) : $signed(_GEN_15575); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15577 = 9'hd8 == cnt[8:0] ? $signed(32'sh3e34) : $signed(_GEN_15576); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15578 = 9'hd9 == cnt[8:0] ? $signed(32'sh3cae) : $signed(_GEN_15577); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15579 = 9'hda == cnt[8:0] ? $signed(32'sh3b27) : $signed(_GEN_15578); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15580 = 9'hdb == cnt[8:0] ? $signed(32'sh399f) : $signed(_GEN_15579); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15581 = 9'hdc == cnt[8:0] ? $signed(32'sh3817) : $signed(_GEN_15580); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15582 = 9'hdd == cnt[8:0] ? $signed(32'sh368e) : $signed(_GEN_15581); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15583 = 9'hde == cnt[8:0] ? $signed(32'sh3505) : $signed(_GEN_15582); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15584 = 9'hdf == cnt[8:0] ? $signed(32'sh337c) : $signed(_GEN_15583); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15585 = 9'he0 == cnt[8:0] ? $signed(32'sh31f1) : $signed(_GEN_15584); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15586 = 9'he1 == cnt[8:0] ? $signed(32'sh3067) : $signed(_GEN_15585); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15587 = 9'he2 == cnt[8:0] ? $signed(32'sh2edc) : $signed(_GEN_15586); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15588 = 9'he3 == cnt[8:0] ? $signed(32'sh2d50) : $signed(_GEN_15587); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15589 = 9'he4 == cnt[8:0] ? $signed(32'sh2bc4) : $signed(_GEN_15588); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15590 = 9'he5 == cnt[8:0] ? $signed(32'sh2a38) : $signed(_GEN_15589); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15591 = 9'he6 == cnt[8:0] ? $signed(32'sh28ab) : $signed(_GEN_15590); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15592 = 9'he7 == cnt[8:0] ? $signed(32'sh271e) : $signed(_GEN_15591); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15593 = 9'he8 == cnt[8:0] ? $signed(32'sh2590) : $signed(_GEN_15592); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15594 = 9'he9 == cnt[8:0] ? $signed(32'sh2402) : $signed(_GEN_15593); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15595 = 9'hea == cnt[8:0] ? $signed(32'sh2274) : $signed(_GEN_15594); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15596 = 9'heb == cnt[8:0] ? $signed(32'sh20e5) : $signed(_GEN_15595); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15597 = 9'hec == cnt[8:0] ? $signed(32'sh1f56) : $signed(_GEN_15596); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15598 = 9'hed == cnt[8:0] ? $signed(32'sh1dc7) : $signed(_GEN_15597); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15599 = 9'hee == cnt[8:0] ? $signed(32'sh1c38) : $signed(_GEN_15598); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15600 = 9'hef == cnt[8:0] ? $signed(32'sh1aa8) : $signed(_GEN_15599); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15601 = 9'hf0 == cnt[8:0] ? $signed(32'sh1918) : $signed(_GEN_15600); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15602 = 9'hf1 == cnt[8:0] ? $signed(32'sh1787) : $signed(_GEN_15601); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15603 = 9'hf2 == cnt[8:0] ? $signed(32'sh15f7) : $signed(_GEN_15602); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15604 = 9'hf3 == cnt[8:0] ? $signed(32'sh1466) : $signed(_GEN_15603); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15605 = 9'hf4 == cnt[8:0] ? $signed(32'sh12d5) : $signed(_GEN_15604); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15606 = 9'hf5 == cnt[8:0] ? $signed(32'sh1144) : $signed(_GEN_15605); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15607 = 9'hf6 == cnt[8:0] ? $signed(32'shfb3) : $signed(_GEN_15606); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15608 = 9'hf7 == cnt[8:0] ? $signed(32'she21) : $signed(_GEN_15607); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15609 = 9'hf8 == cnt[8:0] ? $signed(32'shc90) : $signed(_GEN_15608); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15610 = 9'hf9 == cnt[8:0] ? $signed(32'shafe) : $signed(_GEN_15609); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15611 = 9'hfa == cnt[8:0] ? $signed(32'sh96c) : $signed(_GEN_15610); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15612 = 9'hfb == cnt[8:0] ? $signed(32'sh7da) : $signed(_GEN_15611); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15613 = 9'hfc == cnt[8:0] ? $signed(32'sh648) : $signed(_GEN_15612); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15614 = 9'hfd == cnt[8:0] ? $signed(32'sh4b6) : $signed(_GEN_15613); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15615 = 9'hfe == cnt[8:0] ? $signed(32'sh324) : $signed(_GEN_15614); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15616 = 9'hff == cnt[8:0] ? $signed(32'sh192) : $signed(_GEN_15615); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15617 = 9'h100 == cnt[8:0] ? $signed(32'sh0) : $signed(_GEN_15616); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15618 = 9'h101 == cnt[8:0] ? $signed(-32'sh192) : $signed(_GEN_15617); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15619 = 9'h102 == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_15618); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15620 = 9'h103 == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_15619); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15621 = 9'h104 == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_15620); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15622 = 9'h105 == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_15621); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15623 = 9'h106 == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_15622); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15624 = 9'h107 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_15623); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15625 = 9'h108 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_15624); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15626 = 9'h109 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_15625); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15627 = 9'h10a == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_15626); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15628 = 9'h10b == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_15627); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15629 = 9'h10c == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_15628); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15630 = 9'h10d == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_15629); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15631 = 9'h10e == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_15630); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15632 = 9'h10f == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_15631); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15633 = 9'h110 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_15632); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15634 = 9'h111 == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_15633); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15635 = 9'h112 == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_15634); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15636 = 9'h113 == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_15635); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15637 = 9'h114 == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_15636); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15638 = 9'h115 == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_15637); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15639 = 9'h116 == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_15638); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15640 = 9'h117 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_15639); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15641 = 9'h118 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_15640); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15642 = 9'h119 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_15641); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15643 = 9'h11a == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_15642); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15644 = 9'h11b == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_15643); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15645 = 9'h11c == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_15644); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15646 = 9'h11d == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_15645); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15647 = 9'h11e == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_15646); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15648 = 9'h11f == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_15647); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15649 = 9'h120 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_15648); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15650 = 9'h121 == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_15649); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15651 = 9'h122 == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_15650); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15652 = 9'h123 == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_15651); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15653 = 9'h124 == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_15652); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15654 = 9'h125 == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_15653); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15655 = 9'h126 == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_15654); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15656 = 9'h127 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_15655); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15657 = 9'h128 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_15656); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15658 = 9'h129 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_15657); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15659 = 9'h12a == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_15658); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15660 = 9'h12b == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_15659); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15661 = 9'h12c == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_15660); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15662 = 9'h12d == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_15661); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15663 = 9'h12e == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_15662); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15664 = 9'h12f == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_15663); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15665 = 9'h130 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_15664); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15666 = 9'h131 == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_15665); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15667 = 9'h132 == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_15666); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15668 = 9'h133 == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_15667); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15669 = 9'h134 == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_15668); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15670 = 9'h135 == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_15669); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15671 = 9'h136 == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_15670); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15672 = 9'h137 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_15671); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15673 = 9'h138 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_15672); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15674 = 9'h139 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_15673); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15675 = 9'h13a == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_15674); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15676 = 9'h13b == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_15675); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15677 = 9'h13c == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_15676); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15678 = 9'h13d == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_15677); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15679 = 9'h13e == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_15678); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15680 = 9'h13f == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_15679); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15681 = 9'h140 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_15680); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15682 = 9'h141 == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_15681); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15683 = 9'h142 == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_15682); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15684 = 9'h143 == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_15683); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15685 = 9'h144 == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_15684); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15686 = 9'h145 == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_15685); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15687 = 9'h146 == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_15686); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15688 = 9'h147 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_15687); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15689 = 9'h148 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_15688); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15690 = 9'h149 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_15689); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15691 = 9'h14a == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_15690); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15692 = 9'h14b == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_15691); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15693 = 9'h14c == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_15692); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15694 = 9'h14d == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_15693); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15695 = 9'h14e == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_15694); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15696 = 9'h14f == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_15695); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15697 = 9'h150 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_15696); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15698 = 9'h151 == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_15697); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15699 = 9'h152 == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_15698); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15700 = 9'h153 == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_15699); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15701 = 9'h154 == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_15700); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15702 = 9'h155 == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_15701); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15703 = 9'h156 == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_15702); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15704 = 9'h157 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_15703); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15705 = 9'h158 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_15704); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15706 = 9'h159 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_15705); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15707 = 9'h15a == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_15706); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15708 = 9'h15b == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_15707); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15709 = 9'h15c == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_15708); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15710 = 9'h15d == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_15709); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15711 = 9'h15e == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_15710); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15712 = 9'h15f == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_15711); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15713 = 9'h160 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_15712); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15714 = 9'h161 == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_15713); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15715 = 9'h162 == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_15714); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15716 = 9'h163 == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_15715); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15717 = 9'h164 == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_15716); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15718 = 9'h165 == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_15717); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15719 = 9'h166 == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_15718); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15720 = 9'h167 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_15719); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15721 = 9'h168 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_15720); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15722 = 9'h169 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_15721); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15723 = 9'h16a == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_15722); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15724 = 9'h16b == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_15723); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15725 = 9'h16c == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_15724); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15726 = 9'h16d == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_15725); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15727 = 9'h16e == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_15726); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15728 = 9'h16f == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_15727); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15729 = 9'h170 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_15728); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15730 = 9'h171 == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_15729); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15731 = 9'h172 == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_15730); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15732 = 9'h173 == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_15731); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15733 = 9'h174 == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_15732); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15734 = 9'h175 == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_15733); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15735 = 9'h176 == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_15734); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15736 = 9'h177 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_15735); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15737 = 9'h178 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_15736); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15738 = 9'h179 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_15737); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15739 = 9'h17a == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_15738); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15740 = 9'h17b == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_15739); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15741 = 9'h17c == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_15740); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15742 = 9'h17d == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_15741); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15743 = 9'h17e == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_15742); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15744 = 9'h17f == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_15743); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15745 = 9'h180 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_15744); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15746 = 9'h181 == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_15745); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15747 = 9'h182 == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_15746); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15748 = 9'h183 == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_15747); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15749 = 9'h184 == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_15748); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15750 = 9'h185 == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_15749); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15751 = 9'h186 == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_15750); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15752 = 9'h187 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_15751); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15753 = 9'h188 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_15752); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15754 = 9'h189 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_15753); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15755 = 9'h18a == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_15754); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15756 = 9'h18b == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_15755); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15757 = 9'h18c == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_15756); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15758 = 9'h18d == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_15757); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15759 = 9'h18e == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_15758); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15760 = 9'h18f == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_15759); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15761 = 9'h190 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_15760); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15762 = 9'h191 == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_15761); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15763 = 9'h192 == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_15762); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15764 = 9'h193 == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_15763); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15765 = 9'h194 == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_15764); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15766 = 9'h195 == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_15765); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15767 = 9'h196 == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_15766); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15768 = 9'h197 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_15767); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15769 = 9'h198 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_15768); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15770 = 9'h199 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_15769); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15771 = 9'h19a == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_15770); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15772 = 9'h19b == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_15771); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15773 = 9'h19c == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_15772); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15774 = 9'h19d == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_15773); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15775 = 9'h19e == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_15774); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15776 = 9'h19f == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_15775); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15777 = 9'h1a0 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_15776); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15778 = 9'h1a1 == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_15777); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15779 = 9'h1a2 == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_15778); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15780 = 9'h1a3 == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_15779); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15781 = 9'h1a4 == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_15780); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15782 = 9'h1a5 == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_15781); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15783 = 9'h1a6 == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_15782); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15784 = 9'h1a7 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_15783); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15785 = 9'h1a8 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_15784); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15786 = 9'h1a9 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_15785); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15787 = 9'h1aa == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_15786); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15788 = 9'h1ab == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_15787); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15789 = 9'h1ac == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_15788); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15790 = 9'h1ad == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_15789); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15791 = 9'h1ae == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_15790); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15792 = 9'h1af == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_15791); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15793 = 9'h1b0 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_15792); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15794 = 9'h1b1 == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_15793); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15795 = 9'h1b2 == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_15794); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15796 = 9'h1b3 == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_15795); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15797 = 9'h1b4 == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_15796); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15798 = 9'h1b5 == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_15797); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15799 = 9'h1b6 == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_15798); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15800 = 9'h1b7 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_15799); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15801 = 9'h1b8 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_15800); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15802 = 9'h1b9 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_15801); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15803 = 9'h1ba == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_15802); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15804 = 9'h1bb == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_15803); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15805 = 9'h1bc == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_15804); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15806 = 9'h1bd == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_15805); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15807 = 9'h1be == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_15806); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15808 = 9'h1bf == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_15807); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15809 = 9'h1c0 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_15808); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15810 = 9'h1c1 == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_15809); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15811 = 9'h1c2 == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_15810); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15812 = 9'h1c3 == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_15811); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15813 = 9'h1c4 == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_15812); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15814 = 9'h1c5 == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_15813); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15815 = 9'h1c6 == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_15814); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15816 = 9'h1c7 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_15815); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15817 = 9'h1c8 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_15816); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15818 = 9'h1c9 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_15817); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15819 = 9'h1ca == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_15818); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15820 = 9'h1cb == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_15819); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15821 = 9'h1cc == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_15820); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15822 = 9'h1cd == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_15821); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15823 = 9'h1ce == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_15822); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15824 = 9'h1cf == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_15823); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15825 = 9'h1d0 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_15824); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15826 = 9'h1d1 == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_15825); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15827 = 9'h1d2 == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_15826); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15828 = 9'h1d3 == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_15827); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15829 = 9'h1d4 == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_15828); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15830 = 9'h1d5 == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_15829); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15831 = 9'h1d6 == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_15830); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15832 = 9'h1d7 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_15831); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15833 = 9'h1d8 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_15832); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15834 = 9'h1d9 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_15833); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15835 = 9'h1da == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_15834); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15836 = 9'h1db == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_15835); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15837 = 9'h1dc == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_15836); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15838 = 9'h1dd == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_15837); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15839 = 9'h1de == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_15838); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15840 = 9'h1df == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_15839); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15841 = 9'h1e0 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_15840); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15842 = 9'h1e1 == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_15841); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15843 = 9'h1e2 == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_15842); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15844 = 9'h1e3 == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_15843); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15845 = 9'h1e4 == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_15844); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15846 = 9'h1e5 == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_15845); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15847 = 9'h1e6 == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_15846); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15848 = 9'h1e7 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_15847); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15849 = 9'h1e8 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_15848); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15850 = 9'h1e9 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_15849); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15851 = 9'h1ea == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_15850); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15852 = 9'h1eb == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_15851); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15853 = 9'h1ec == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_15852); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15854 = 9'h1ed == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_15853); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15855 = 9'h1ee == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_15854); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15856 = 9'h1ef == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_15855); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15857 = 9'h1f0 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_15856); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15858 = 9'h1f1 == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_15857); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15859 = 9'h1f2 == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_15858); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15860 = 9'h1f3 == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_15859); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15861 = 9'h1f4 == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_15860); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15862 = 9'h1f5 == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_15861); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15863 = 9'h1f6 == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_15862); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15864 = 9'h1f7 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_15863); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15865 = 9'h1f8 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_15864); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15866 = 9'h1f9 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_15865); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15867 = 9'h1fa == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_15866); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15868 = 9'h1fb == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_15867); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15869 = 9'h1fc == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_15868); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15870 = 9'h1fd == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_15869); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15871 = 9'h1fe == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_15870); // @[FFT.scala 34:12]
  wire [31:0] _GEN_15874 = 9'h1 == cnt[8:0] ? $signed(-32'sh192) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15875 = 9'h2 == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_15874); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15876 = 9'h3 == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_15875); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15877 = 9'h4 == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_15876); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15878 = 9'h5 == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_15877); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15879 = 9'h6 == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_15878); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15880 = 9'h7 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_15879); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15881 = 9'h8 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_15880); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15882 = 9'h9 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_15881); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15883 = 9'ha == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_15882); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15884 = 9'hb == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_15883); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15885 = 9'hc == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_15884); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15886 = 9'hd == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_15885); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15887 = 9'he == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_15886); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15888 = 9'hf == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_15887); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15889 = 9'h10 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_15888); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15890 = 9'h11 == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_15889); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15891 = 9'h12 == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_15890); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15892 = 9'h13 == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_15891); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15893 = 9'h14 == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_15892); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15894 = 9'h15 == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_15893); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15895 = 9'h16 == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_15894); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15896 = 9'h17 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_15895); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15897 = 9'h18 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_15896); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15898 = 9'h19 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_15897); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15899 = 9'h1a == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_15898); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15900 = 9'h1b == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_15899); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15901 = 9'h1c == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_15900); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15902 = 9'h1d == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_15901); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15903 = 9'h1e == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_15902); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15904 = 9'h1f == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_15903); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15905 = 9'h20 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_15904); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15906 = 9'h21 == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_15905); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15907 = 9'h22 == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_15906); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15908 = 9'h23 == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_15907); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15909 = 9'h24 == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_15908); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15910 = 9'h25 == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_15909); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15911 = 9'h26 == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_15910); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15912 = 9'h27 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_15911); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15913 = 9'h28 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_15912); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15914 = 9'h29 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_15913); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15915 = 9'h2a == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_15914); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15916 = 9'h2b == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_15915); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15917 = 9'h2c == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_15916); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15918 = 9'h2d == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_15917); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15919 = 9'h2e == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_15918); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15920 = 9'h2f == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_15919); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15921 = 9'h30 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_15920); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15922 = 9'h31 == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_15921); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15923 = 9'h32 == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_15922); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15924 = 9'h33 == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_15923); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15925 = 9'h34 == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_15924); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15926 = 9'h35 == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_15925); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15927 = 9'h36 == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_15926); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15928 = 9'h37 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_15927); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15929 = 9'h38 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_15928); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15930 = 9'h39 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_15929); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15931 = 9'h3a == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_15930); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15932 = 9'h3b == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_15931); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15933 = 9'h3c == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_15932); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15934 = 9'h3d == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_15933); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15935 = 9'h3e == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_15934); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15936 = 9'h3f == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_15935); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15937 = 9'h40 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_15936); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15938 = 9'h41 == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_15937); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15939 = 9'h42 == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_15938); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15940 = 9'h43 == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_15939); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15941 = 9'h44 == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_15940); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15942 = 9'h45 == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_15941); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15943 = 9'h46 == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_15942); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15944 = 9'h47 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_15943); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15945 = 9'h48 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_15944); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15946 = 9'h49 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_15945); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15947 = 9'h4a == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_15946); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15948 = 9'h4b == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_15947); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15949 = 9'h4c == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_15948); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15950 = 9'h4d == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_15949); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15951 = 9'h4e == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_15950); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15952 = 9'h4f == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_15951); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15953 = 9'h50 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_15952); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15954 = 9'h51 == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_15953); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15955 = 9'h52 == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_15954); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15956 = 9'h53 == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_15955); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15957 = 9'h54 == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_15956); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15958 = 9'h55 == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_15957); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15959 = 9'h56 == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_15958); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15960 = 9'h57 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_15959); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15961 = 9'h58 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_15960); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15962 = 9'h59 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_15961); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15963 = 9'h5a == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_15962); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15964 = 9'h5b == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_15963); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15965 = 9'h5c == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_15964); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15966 = 9'h5d == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_15965); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15967 = 9'h5e == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_15966); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15968 = 9'h5f == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_15967); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15969 = 9'h60 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_15968); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15970 = 9'h61 == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_15969); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15971 = 9'h62 == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_15970); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15972 = 9'h63 == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_15971); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15973 = 9'h64 == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_15972); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15974 = 9'h65 == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_15973); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15975 = 9'h66 == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_15974); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15976 = 9'h67 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_15975); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15977 = 9'h68 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_15976); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15978 = 9'h69 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_15977); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15979 = 9'h6a == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_15978); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15980 = 9'h6b == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_15979); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15981 = 9'h6c == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_15980); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15982 = 9'h6d == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_15981); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15983 = 9'h6e == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_15982); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15984 = 9'h6f == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_15983); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15985 = 9'h70 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_15984); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15986 = 9'h71 == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_15985); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15987 = 9'h72 == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_15986); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15988 = 9'h73 == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_15987); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15989 = 9'h74 == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_15988); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15990 = 9'h75 == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_15989); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15991 = 9'h76 == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_15990); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15992 = 9'h77 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_15991); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15993 = 9'h78 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_15992); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15994 = 9'h79 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_15993); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15995 = 9'h7a == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_15994); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15996 = 9'h7b == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_15995); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15997 = 9'h7c == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_15996); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15998 = 9'h7d == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_15997); // @[FFT.scala 35:12]
  wire [31:0] _GEN_15999 = 9'h7e == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_15998); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16000 = 9'h7f == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_15999); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16001 = 9'h80 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_16000); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16002 = 9'h81 == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_16001); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16003 = 9'h82 == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_16002); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16004 = 9'h83 == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_16003); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16005 = 9'h84 == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_16004); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16006 = 9'h85 == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_16005); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16007 = 9'h86 == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_16006); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16008 = 9'h87 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_16007); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16009 = 9'h88 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_16008); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16010 = 9'h89 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_16009); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16011 = 9'h8a == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_16010); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16012 = 9'h8b == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_16011); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16013 = 9'h8c == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_16012); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16014 = 9'h8d == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_16013); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16015 = 9'h8e == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_16014); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16016 = 9'h8f == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_16015); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16017 = 9'h90 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_16016); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16018 = 9'h91 == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_16017); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16019 = 9'h92 == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_16018); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16020 = 9'h93 == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_16019); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16021 = 9'h94 == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_16020); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16022 = 9'h95 == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_16021); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16023 = 9'h96 == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_16022); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16024 = 9'h97 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_16023); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16025 = 9'h98 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_16024); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16026 = 9'h99 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_16025); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16027 = 9'h9a == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_16026); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16028 = 9'h9b == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_16027); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16029 = 9'h9c == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_16028); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16030 = 9'h9d == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_16029); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16031 = 9'h9e == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_16030); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16032 = 9'h9f == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_16031); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16033 = 9'ha0 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_16032); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16034 = 9'ha1 == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_16033); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16035 = 9'ha2 == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_16034); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16036 = 9'ha3 == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_16035); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16037 = 9'ha4 == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_16036); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16038 = 9'ha5 == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_16037); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16039 = 9'ha6 == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_16038); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16040 = 9'ha7 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_16039); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16041 = 9'ha8 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_16040); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16042 = 9'ha9 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_16041); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16043 = 9'haa == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_16042); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16044 = 9'hab == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_16043); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16045 = 9'hac == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_16044); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16046 = 9'had == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_16045); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16047 = 9'hae == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_16046); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16048 = 9'haf == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_16047); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16049 = 9'hb0 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_16048); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16050 = 9'hb1 == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_16049); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16051 = 9'hb2 == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_16050); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16052 = 9'hb3 == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_16051); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16053 = 9'hb4 == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_16052); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16054 = 9'hb5 == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_16053); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16055 = 9'hb6 == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_16054); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16056 = 9'hb7 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_16055); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16057 = 9'hb8 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_16056); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16058 = 9'hb9 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_16057); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16059 = 9'hba == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_16058); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16060 = 9'hbb == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_16059); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16061 = 9'hbc == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_16060); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16062 = 9'hbd == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_16061); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16063 = 9'hbe == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_16062); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16064 = 9'hbf == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_16063); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16065 = 9'hc0 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_16064); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16066 = 9'hc1 == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_16065); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16067 = 9'hc2 == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_16066); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16068 = 9'hc3 == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_16067); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16069 = 9'hc4 == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_16068); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16070 = 9'hc5 == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_16069); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16071 = 9'hc6 == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_16070); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16072 = 9'hc7 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_16071); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16073 = 9'hc8 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_16072); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16074 = 9'hc9 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_16073); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16075 = 9'hca == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_16074); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16076 = 9'hcb == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_16075); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16077 = 9'hcc == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_16076); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16078 = 9'hcd == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_16077); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16079 = 9'hce == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_16078); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16080 = 9'hcf == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_16079); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16081 = 9'hd0 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_16080); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16082 = 9'hd1 == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_16081); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16083 = 9'hd2 == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_16082); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16084 = 9'hd3 == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_16083); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16085 = 9'hd4 == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_16084); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16086 = 9'hd5 == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_16085); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16087 = 9'hd6 == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_16086); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16088 = 9'hd7 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_16087); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16089 = 9'hd8 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_16088); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16090 = 9'hd9 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_16089); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16091 = 9'hda == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_16090); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16092 = 9'hdb == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_16091); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16093 = 9'hdc == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_16092); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16094 = 9'hdd == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_16093); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16095 = 9'hde == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_16094); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16096 = 9'hdf == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_16095); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16097 = 9'he0 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_16096); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16098 = 9'he1 == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_16097); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16099 = 9'he2 == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_16098); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16100 = 9'he3 == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_16099); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16101 = 9'he4 == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_16100); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16102 = 9'he5 == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_16101); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16103 = 9'he6 == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_16102); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16104 = 9'he7 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_16103); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16105 = 9'he8 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_16104); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16106 = 9'he9 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_16105); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16107 = 9'hea == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_16106); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16108 = 9'heb == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_16107); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16109 = 9'hec == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_16108); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16110 = 9'hed == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_16109); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16111 = 9'hee == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_16110); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16112 = 9'hef == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_16111); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16113 = 9'hf0 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_16112); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16114 = 9'hf1 == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_16113); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16115 = 9'hf2 == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_16114); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16116 = 9'hf3 == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_16115); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16117 = 9'hf4 == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_16116); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16118 = 9'hf5 == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_16117); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16119 = 9'hf6 == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_16118); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16120 = 9'hf7 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_16119); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16121 = 9'hf8 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_16120); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16122 = 9'hf9 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_16121); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16123 = 9'hfa == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_16122); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16124 = 9'hfb == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_16123); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16125 = 9'hfc == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_16124); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16126 = 9'hfd == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_16125); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16127 = 9'hfe == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_16126); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16128 = 9'hff == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_16127); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16129 = 9'h100 == cnt[8:0] ? $signed(-32'sh10000) : $signed(_GEN_16128); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16130 = 9'h101 == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_16129); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16131 = 9'h102 == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_16130); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16132 = 9'h103 == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_16131); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16133 = 9'h104 == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_16132); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16134 = 9'h105 == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_16133); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16135 = 9'h106 == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_16134); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16136 = 9'h107 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_16135); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16137 = 9'h108 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_16136); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16138 = 9'h109 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_16137); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16139 = 9'h10a == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_16138); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16140 = 9'h10b == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_16139); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16141 = 9'h10c == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_16140); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16142 = 9'h10d == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_16141); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16143 = 9'h10e == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_16142); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16144 = 9'h10f == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_16143); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16145 = 9'h110 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_16144); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16146 = 9'h111 == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_16145); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16147 = 9'h112 == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_16146); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16148 = 9'h113 == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_16147); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16149 = 9'h114 == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_16148); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16150 = 9'h115 == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_16149); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16151 = 9'h116 == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_16150); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16152 = 9'h117 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_16151); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16153 = 9'h118 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_16152); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16154 = 9'h119 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_16153); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16155 = 9'h11a == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_16154); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16156 = 9'h11b == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_16155); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16157 = 9'h11c == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_16156); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16158 = 9'h11d == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_16157); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16159 = 9'h11e == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_16158); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16160 = 9'h11f == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_16159); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16161 = 9'h120 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_16160); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16162 = 9'h121 == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_16161); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16163 = 9'h122 == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_16162); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16164 = 9'h123 == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_16163); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16165 = 9'h124 == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_16164); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16166 = 9'h125 == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_16165); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16167 = 9'h126 == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_16166); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16168 = 9'h127 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_16167); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16169 = 9'h128 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_16168); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16170 = 9'h129 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_16169); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16171 = 9'h12a == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_16170); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16172 = 9'h12b == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_16171); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16173 = 9'h12c == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_16172); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16174 = 9'h12d == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_16173); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16175 = 9'h12e == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_16174); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16176 = 9'h12f == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_16175); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16177 = 9'h130 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_16176); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16178 = 9'h131 == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_16177); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16179 = 9'h132 == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_16178); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16180 = 9'h133 == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_16179); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16181 = 9'h134 == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_16180); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16182 = 9'h135 == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_16181); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16183 = 9'h136 == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_16182); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16184 = 9'h137 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_16183); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16185 = 9'h138 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_16184); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16186 = 9'h139 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_16185); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16187 = 9'h13a == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_16186); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16188 = 9'h13b == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_16187); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16189 = 9'h13c == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_16188); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16190 = 9'h13d == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_16189); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16191 = 9'h13e == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_16190); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16192 = 9'h13f == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_16191); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16193 = 9'h140 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_16192); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16194 = 9'h141 == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_16193); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16195 = 9'h142 == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_16194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16196 = 9'h143 == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_16195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16197 = 9'h144 == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_16196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16198 = 9'h145 == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_16197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16199 = 9'h146 == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_16198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16200 = 9'h147 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_16199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16201 = 9'h148 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_16200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16202 = 9'h149 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_16201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16203 = 9'h14a == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_16202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16204 = 9'h14b == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_16203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16205 = 9'h14c == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_16204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16206 = 9'h14d == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_16205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16207 = 9'h14e == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_16206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16208 = 9'h14f == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_16207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16209 = 9'h150 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_16208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16210 = 9'h151 == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_16209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16211 = 9'h152 == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_16210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16212 = 9'h153 == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_16211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16213 = 9'h154 == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_16212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16214 = 9'h155 == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_16213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16215 = 9'h156 == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_16214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16216 = 9'h157 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_16215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16217 = 9'h158 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_16216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16218 = 9'h159 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_16217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16219 = 9'h15a == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_16218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16220 = 9'h15b == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_16219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16221 = 9'h15c == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_16220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16222 = 9'h15d == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_16221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16223 = 9'h15e == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_16222); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16224 = 9'h15f == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_16223); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16225 = 9'h160 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_16224); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16226 = 9'h161 == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_16225); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16227 = 9'h162 == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_16226); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16228 = 9'h163 == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_16227); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16229 = 9'h164 == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_16228); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16230 = 9'h165 == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_16229); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16231 = 9'h166 == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_16230); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16232 = 9'h167 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_16231); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16233 = 9'h168 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_16232); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16234 = 9'h169 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_16233); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16235 = 9'h16a == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_16234); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16236 = 9'h16b == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_16235); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16237 = 9'h16c == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_16236); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16238 = 9'h16d == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_16237); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16239 = 9'h16e == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_16238); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16240 = 9'h16f == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_16239); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16241 = 9'h170 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_16240); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16242 = 9'h171 == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_16241); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16243 = 9'h172 == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_16242); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16244 = 9'h173 == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_16243); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16245 = 9'h174 == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_16244); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16246 = 9'h175 == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_16245); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16247 = 9'h176 == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_16246); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16248 = 9'h177 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_16247); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16249 = 9'h178 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_16248); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16250 = 9'h179 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_16249); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16251 = 9'h17a == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_16250); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16252 = 9'h17b == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_16251); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16253 = 9'h17c == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_16252); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16254 = 9'h17d == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_16253); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16255 = 9'h17e == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_16254); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16256 = 9'h17f == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_16255); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16257 = 9'h180 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_16256); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16258 = 9'h181 == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_16257); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16259 = 9'h182 == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_16258); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16260 = 9'h183 == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_16259); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16261 = 9'h184 == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_16260); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16262 = 9'h185 == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_16261); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16263 = 9'h186 == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_16262); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16264 = 9'h187 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_16263); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16265 = 9'h188 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_16264); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16266 = 9'h189 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_16265); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16267 = 9'h18a == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_16266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16268 = 9'h18b == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_16267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16269 = 9'h18c == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_16268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16270 = 9'h18d == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_16269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16271 = 9'h18e == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_16270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16272 = 9'h18f == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_16271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16273 = 9'h190 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_16272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16274 = 9'h191 == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_16273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16275 = 9'h192 == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_16274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16276 = 9'h193 == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_16275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16277 = 9'h194 == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_16276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16278 = 9'h195 == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_16277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16279 = 9'h196 == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_16278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16280 = 9'h197 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_16279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16281 = 9'h198 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_16280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16282 = 9'h199 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_16281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16283 = 9'h19a == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_16282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16284 = 9'h19b == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_16283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16285 = 9'h19c == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_16284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16286 = 9'h19d == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_16285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16287 = 9'h19e == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_16286); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16288 = 9'h19f == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_16287); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16289 = 9'h1a0 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_16288); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16290 = 9'h1a1 == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_16289); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16291 = 9'h1a2 == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_16290); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16292 = 9'h1a3 == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_16291); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16293 = 9'h1a4 == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_16292); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16294 = 9'h1a5 == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_16293); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16295 = 9'h1a6 == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_16294); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16296 = 9'h1a7 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_16295); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16297 = 9'h1a8 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_16296); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16298 = 9'h1a9 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_16297); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16299 = 9'h1aa == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_16298); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16300 = 9'h1ab == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_16299); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16301 = 9'h1ac == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_16300); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16302 = 9'h1ad == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_16301); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16303 = 9'h1ae == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_16302); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16304 = 9'h1af == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_16303); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16305 = 9'h1b0 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_16304); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16306 = 9'h1b1 == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_16305); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16307 = 9'h1b2 == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_16306); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16308 = 9'h1b3 == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_16307); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16309 = 9'h1b4 == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_16308); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16310 = 9'h1b5 == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_16309); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16311 = 9'h1b6 == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_16310); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16312 = 9'h1b7 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_16311); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16313 = 9'h1b8 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_16312); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16314 = 9'h1b9 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_16313); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16315 = 9'h1ba == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_16314); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16316 = 9'h1bb == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_16315); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16317 = 9'h1bc == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_16316); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16318 = 9'h1bd == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_16317); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16319 = 9'h1be == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_16318); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16320 = 9'h1bf == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_16319); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16321 = 9'h1c0 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_16320); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16322 = 9'h1c1 == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_16321); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16323 = 9'h1c2 == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_16322); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16324 = 9'h1c3 == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_16323); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16325 = 9'h1c4 == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_16324); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16326 = 9'h1c5 == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_16325); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16327 = 9'h1c6 == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_16326); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16328 = 9'h1c7 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_16327); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16329 = 9'h1c8 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_16328); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16330 = 9'h1c9 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_16329); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16331 = 9'h1ca == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_16330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16332 = 9'h1cb == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_16331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16333 = 9'h1cc == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_16332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16334 = 9'h1cd == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_16333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16335 = 9'h1ce == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_16334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16336 = 9'h1cf == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_16335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16337 = 9'h1d0 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_16336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16338 = 9'h1d1 == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_16337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16339 = 9'h1d2 == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_16338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16340 = 9'h1d3 == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_16339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16341 = 9'h1d4 == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_16340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16342 = 9'h1d5 == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_16341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16343 = 9'h1d6 == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_16342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16344 = 9'h1d7 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_16343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16345 = 9'h1d8 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_16344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16346 = 9'h1d9 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_16345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16347 = 9'h1da == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_16346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16348 = 9'h1db == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_16347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16349 = 9'h1dc == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_16348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16350 = 9'h1dd == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_16349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16351 = 9'h1de == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_16350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16352 = 9'h1df == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_16351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16353 = 9'h1e0 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_16352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16354 = 9'h1e1 == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_16353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16355 = 9'h1e2 == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_16354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16356 = 9'h1e3 == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_16355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16357 = 9'h1e4 == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_16356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16358 = 9'h1e5 == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_16357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16359 = 9'h1e6 == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_16358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16360 = 9'h1e7 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_16359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16361 = 9'h1e8 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_16360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16362 = 9'h1e9 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_16361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16363 = 9'h1ea == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_16362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16364 = 9'h1eb == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_16363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16365 = 9'h1ec == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_16364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16366 = 9'h1ed == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_16365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16367 = 9'h1ee == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_16366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16368 = 9'h1ef == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_16367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16369 = 9'h1f0 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_16368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16370 = 9'h1f1 == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_16369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16371 = 9'h1f2 == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_16370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16372 = 9'h1f3 == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_16371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16373 = 9'h1f4 == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_16372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16374 = 9'h1f5 == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_16373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16375 = 9'h1f6 == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_16374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16376 = 9'h1f7 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_16375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16377 = 9'h1f8 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_16376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16378 = 9'h1f9 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_16377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16379 = 9'h1fa == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_16378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16380 = 9'h1fb == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_16379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16381 = 9'h1fc == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_16380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16382 = 9'h1fd == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_16381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_16383 = 9'h1fe == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_16382); // @[FFT.scala 35:12]
  reg [31:0] _T_4811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9218;
  reg [31:0] _T_4811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9219;
  reg [31:0] _T_4812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9220;
  reg [31:0] _T_4812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9221;
  reg [31:0] _T_4813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9222;
  reg [31:0] _T_4813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9223;
  reg [31:0] _T_4814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9224;
  reg [31:0] _T_4814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9225;
  reg [31:0] _T_4815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9226;
  reg [31:0] _T_4815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9227;
  reg [31:0] _T_4816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9228;
  reg [31:0] _T_4816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9229;
  reg [31:0] _T_4817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9230;
  reg [31:0] _T_4817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9231;
  reg [31:0] _T_4818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9232;
  reg [31:0] _T_4818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9233;
  reg [31:0] _T_4819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9234;
  reg [31:0] _T_4819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9235;
  reg [31:0] _T_4820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9236;
  reg [31:0] _T_4820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9237;
  reg [31:0] _T_4821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9238;
  reg [31:0] _T_4821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9239;
  reg [31:0] _T_4822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9240;
  reg [31:0] _T_4822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9241;
  reg [31:0] _T_4823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9242;
  reg [31:0] _T_4823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9243;
  reg [31:0] _T_4824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9244;
  reg [31:0] _T_4824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9245;
  reg [31:0] _T_4825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9246;
  reg [31:0] _T_4825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9247;
  reg [31:0] _T_4826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9248;
  reg [31:0] _T_4826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9249;
  reg [31:0] _T_4827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9250;
  reg [31:0] _T_4827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9251;
  reg [31:0] _T_4828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9252;
  reg [31:0] _T_4828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9253;
  reg [31:0] _T_4829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9254;
  reg [31:0] _T_4829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9255;
  reg [31:0] _T_4830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9256;
  reg [31:0] _T_4830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9257;
  reg [31:0] _T_4831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9258;
  reg [31:0] _T_4831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9259;
  reg [31:0] _T_4832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9260;
  reg [31:0] _T_4832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9261;
  reg [31:0] _T_4833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9262;
  reg [31:0] _T_4833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9263;
  reg [31:0] _T_4834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9264;
  reg [31:0] _T_4834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9265;
  reg [31:0] _T_4835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9266;
  reg [31:0] _T_4835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9267;
  reg [31:0] _T_4836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9268;
  reg [31:0] _T_4836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9269;
  reg [31:0] _T_4837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9270;
  reg [31:0] _T_4837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9271;
  reg [31:0] _T_4838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9272;
  reg [31:0] _T_4838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9273;
  reg [31:0] _T_4839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9274;
  reg [31:0] _T_4839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9275;
  reg [31:0] _T_4840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9276;
  reg [31:0] _T_4840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9277;
  reg [31:0] _T_4841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9278;
  reg [31:0] _T_4841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9279;
  reg [31:0] _T_4842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9280;
  reg [31:0] _T_4842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9281;
  reg [31:0] _T_4843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9282;
  reg [31:0] _T_4843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9283;
  reg [31:0] _T_4844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9284;
  reg [31:0] _T_4844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9285;
  reg [31:0] _T_4845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9286;
  reg [31:0] _T_4845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9287;
  reg [31:0] _T_4846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9288;
  reg [31:0] _T_4846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9289;
  reg [31:0] _T_4847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9290;
  reg [31:0] _T_4847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9291;
  reg [31:0] _T_4848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9292;
  reg [31:0] _T_4848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9293;
  reg [31:0] _T_4849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9294;
  reg [31:0] _T_4849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9295;
  reg [31:0] _T_4850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9296;
  reg [31:0] _T_4850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9297;
  reg [31:0] _T_4851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9298;
  reg [31:0] _T_4851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9299;
  reg [31:0] _T_4852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9300;
  reg [31:0] _T_4852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9301;
  reg [31:0] _T_4853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9302;
  reg [31:0] _T_4853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9303;
  reg [31:0] _T_4854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9304;
  reg [31:0] _T_4854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9305;
  reg [31:0] _T_4855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9306;
  reg [31:0] _T_4855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9307;
  reg [31:0] _T_4856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9308;
  reg [31:0] _T_4856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9309;
  reg [31:0] _T_4857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9310;
  reg [31:0] _T_4857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9311;
  reg [31:0] _T_4858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9312;
  reg [31:0] _T_4858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9313;
  reg [31:0] _T_4859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9314;
  reg [31:0] _T_4859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9315;
  reg [31:0] _T_4860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9316;
  reg [31:0] _T_4860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9317;
  reg [31:0] _T_4861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9318;
  reg [31:0] _T_4861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9319;
  reg [31:0] _T_4862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9320;
  reg [31:0] _T_4862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9321;
  reg [31:0] _T_4863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9322;
  reg [31:0] _T_4863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9323;
  reg [31:0] _T_4864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9324;
  reg [31:0] _T_4864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9325;
  reg [31:0] _T_4865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9326;
  reg [31:0] _T_4865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9327;
  reg [31:0] _T_4866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9328;
  reg [31:0] _T_4866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9329;
  reg [31:0] _T_4867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9330;
  reg [31:0] _T_4867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9331;
  reg [31:0] _T_4868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9332;
  reg [31:0] _T_4868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9333;
  reg [31:0] _T_4869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9334;
  reg [31:0] _T_4869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9335;
  reg [31:0] _T_4870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9336;
  reg [31:0] _T_4870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9337;
  reg [31:0] _T_4871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9338;
  reg [31:0] _T_4871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9339;
  reg [31:0] _T_4872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9340;
  reg [31:0] _T_4872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9341;
  reg [31:0] _T_4873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9342;
  reg [31:0] _T_4873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9343;
  reg [31:0] _T_4874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9344;
  reg [31:0] _T_4874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9345;
  reg [31:0] _T_4875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9346;
  reg [31:0] _T_4875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9347;
  reg [31:0] _T_4876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9348;
  reg [31:0] _T_4876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9349;
  reg [31:0] _T_4877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9350;
  reg [31:0] _T_4877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9351;
  reg [31:0] _T_4878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9352;
  reg [31:0] _T_4878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9353;
  reg [31:0] _T_4879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9354;
  reg [31:0] _T_4879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9355;
  reg [31:0] _T_4880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9356;
  reg [31:0] _T_4880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9357;
  reg [31:0] _T_4881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9358;
  reg [31:0] _T_4881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9359;
  reg [31:0] _T_4882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9360;
  reg [31:0] _T_4882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9361;
  reg [31:0] _T_4883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9362;
  reg [31:0] _T_4883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9363;
  reg [31:0] _T_4884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9364;
  reg [31:0] _T_4884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9365;
  reg [31:0] _T_4885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9366;
  reg [31:0] _T_4885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9367;
  reg [31:0] _T_4886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9368;
  reg [31:0] _T_4886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9369;
  reg [31:0] _T_4887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9370;
  reg [31:0] _T_4887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9371;
  reg [31:0] _T_4888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9372;
  reg [31:0] _T_4888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9373;
  reg [31:0] _T_4889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9374;
  reg [31:0] _T_4889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9375;
  reg [31:0] _T_4890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9376;
  reg [31:0] _T_4890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9377;
  reg [31:0] _T_4891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9378;
  reg [31:0] _T_4891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9379;
  reg [31:0] _T_4892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9380;
  reg [31:0] _T_4892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9381;
  reg [31:0] _T_4893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9382;
  reg [31:0] _T_4893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9383;
  reg [31:0] _T_4894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9384;
  reg [31:0] _T_4894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9385;
  reg [31:0] _T_4895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9386;
  reg [31:0] _T_4895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9387;
  reg [31:0] _T_4896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9388;
  reg [31:0] _T_4896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9389;
  reg [31:0] _T_4897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9390;
  reg [31:0] _T_4897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9391;
  reg [31:0] _T_4898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9392;
  reg [31:0] _T_4898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9393;
  reg [31:0] _T_4899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9394;
  reg [31:0] _T_4899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9395;
  reg [31:0] _T_4900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9396;
  reg [31:0] _T_4900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9397;
  reg [31:0] _T_4901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9398;
  reg [31:0] _T_4901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9399;
  reg [31:0] _T_4902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9400;
  reg [31:0] _T_4902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9401;
  reg [31:0] _T_4903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9402;
  reg [31:0] _T_4903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9403;
  reg [31:0] _T_4904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9404;
  reg [31:0] _T_4904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9405;
  reg [31:0] _T_4905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9406;
  reg [31:0] _T_4905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9407;
  reg [31:0] _T_4906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9408;
  reg [31:0] _T_4906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9409;
  reg [31:0] _T_4907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9410;
  reg [31:0] _T_4907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9411;
  reg [31:0] _T_4908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9412;
  reg [31:0] _T_4908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9413;
  reg [31:0] _T_4909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9414;
  reg [31:0] _T_4909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9415;
  reg [31:0] _T_4910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9416;
  reg [31:0] _T_4910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9417;
  reg [31:0] _T_4911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9418;
  reg [31:0] _T_4911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9419;
  reg [31:0] _T_4912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9420;
  reg [31:0] _T_4912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9421;
  reg [31:0] _T_4913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9422;
  reg [31:0] _T_4913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9423;
  reg [31:0] _T_4914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9424;
  reg [31:0] _T_4914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9425;
  reg [31:0] _T_4915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9426;
  reg [31:0] _T_4915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9427;
  reg [31:0] _T_4916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9428;
  reg [31:0] _T_4916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9429;
  reg [31:0] _T_4917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9430;
  reg [31:0] _T_4917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9431;
  reg [31:0] _T_4918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9432;
  reg [31:0] _T_4918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9433;
  reg [31:0] _T_4919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9434;
  reg [31:0] _T_4919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9435;
  reg [31:0] _T_4920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9436;
  reg [31:0] _T_4920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9437;
  reg [31:0] _T_4921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9438;
  reg [31:0] _T_4921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9439;
  reg [31:0] _T_4922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9440;
  reg [31:0] _T_4922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9441;
  reg [31:0] _T_4923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9442;
  reg [31:0] _T_4923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9443;
  reg [31:0] _T_4924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9444;
  reg [31:0] _T_4924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9445;
  reg [31:0] _T_4925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9446;
  reg [31:0] _T_4925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9447;
  reg [31:0] _T_4926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9448;
  reg [31:0] _T_4926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9449;
  reg [31:0] _T_4927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9450;
  reg [31:0] _T_4927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9451;
  reg [31:0] _T_4928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9452;
  reg [31:0] _T_4928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9453;
  reg [31:0] _T_4929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9454;
  reg [31:0] _T_4929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9455;
  reg [31:0] _T_4930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9456;
  reg [31:0] _T_4930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9457;
  reg [31:0] _T_4931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9458;
  reg [31:0] _T_4931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9459;
  reg [31:0] _T_4932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9460;
  reg [31:0] _T_4932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9461;
  reg [31:0] _T_4933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9462;
  reg [31:0] _T_4933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9463;
  reg [31:0] _T_4934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9464;
  reg [31:0] _T_4934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9465;
  reg [31:0] _T_4935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9466;
  reg [31:0] _T_4935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9467;
  reg [31:0] _T_4936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9468;
  reg [31:0] _T_4936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9469;
  reg [31:0] _T_4937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9470;
  reg [31:0] _T_4937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9471;
  reg [31:0] _T_4938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9472;
  reg [31:0] _T_4938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9473;
  reg [31:0] _T_4939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9474;
  reg [31:0] _T_4939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9475;
  reg [31:0] _T_4940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9476;
  reg [31:0] _T_4940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9477;
  reg [31:0] _T_4941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9478;
  reg [31:0] _T_4941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9479;
  reg [31:0] _T_4942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9480;
  reg [31:0] _T_4942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9481;
  reg [31:0] _T_4943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9482;
  reg [31:0] _T_4943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9483;
  reg [31:0] _T_4944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9484;
  reg [31:0] _T_4944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9485;
  reg [31:0] _T_4945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9486;
  reg [31:0] _T_4945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9487;
  reg [31:0] _T_4946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9488;
  reg [31:0] _T_4946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9489;
  reg [31:0] _T_4947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9490;
  reg [31:0] _T_4947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9491;
  reg [31:0] _T_4948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9492;
  reg [31:0] _T_4948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9493;
  reg [31:0] _T_4949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9494;
  reg [31:0] _T_4949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9495;
  reg [31:0] _T_4950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9496;
  reg [31:0] _T_4950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9497;
  reg [31:0] _T_4951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9498;
  reg [31:0] _T_4951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9499;
  reg [31:0] _T_4952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9500;
  reg [31:0] _T_4952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9501;
  reg [31:0] _T_4953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9502;
  reg [31:0] _T_4953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9503;
  reg [31:0] _T_4954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9504;
  reg [31:0] _T_4954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9505;
  reg [31:0] _T_4955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9506;
  reg [31:0] _T_4955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9507;
  reg [31:0] _T_4956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9508;
  reg [31:0] _T_4956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9509;
  reg [31:0] _T_4957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9510;
  reg [31:0] _T_4957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9511;
  reg [31:0] _T_4958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9512;
  reg [31:0] _T_4958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9513;
  reg [31:0] _T_4959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9514;
  reg [31:0] _T_4959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9515;
  reg [31:0] _T_4960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9516;
  reg [31:0] _T_4960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9517;
  reg [31:0] _T_4961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9518;
  reg [31:0] _T_4961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9519;
  reg [31:0] _T_4962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9520;
  reg [31:0] _T_4962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9521;
  reg [31:0] _T_4963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9522;
  reg [31:0] _T_4963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9523;
  reg [31:0] _T_4964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9524;
  reg [31:0] _T_4964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9525;
  reg [31:0] _T_4965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9526;
  reg [31:0] _T_4965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9527;
  reg [31:0] _T_4966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9528;
  reg [31:0] _T_4966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9529;
  reg [31:0] _T_4967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9530;
  reg [31:0] _T_4967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9531;
  reg [31:0] _T_4968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9532;
  reg [31:0] _T_4968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9533;
  reg [31:0] _T_4969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9534;
  reg [31:0] _T_4969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9535;
  reg [31:0] _T_4970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9536;
  reg [31:0] _T_4970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9537;
  reg [31:0] _T_4971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9538;
  reg [31:0] _T_4971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9539;
  reg [31:0] _T_4972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9540;
  reg [31:0] _T_4972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9541;
  reg [31:0] _T_4973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9542;
  reg [31:0] _T_4973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9543;
  reg [31:0] _T_4974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9544;
  reg [31:0] _T_4974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9545;
  reg [31:0] _T_4975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9546;
  reg [31:0] _T_4975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9547;
  reg [31:0] _T_4976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9548;
  reg [31:0] _T_4976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9549;
  reg [31:0] _T_4977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9550;
  reg [31:0] _T_4977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9551;
  reg [31:0] _T_4978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9552;
  reg [31:0] _T_4978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9553;
  reg [31:0] _T_4979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9554;
  reg [31:0] _T_4979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9555;
  reg [31:0] _T_4980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9556;
  reg [31:0] _T_4980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9557;
  reg [31:0] _T_4981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9558;
  reg [31:0] _T_4981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9559;
  reg [31:0] _T_4982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9560;
  reg [31:0] _T_4982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9561;
  reg [31:0] _T_4983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9562;
  reg [31:0] _T_4983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9563;
  reg [31:0] _T_4984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9564;
  reg [31:0] _T_4984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9565;
  reg [31:0] _T_4985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9566;
  reg [31:0] _T_4985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9567;
  reg [31:0] _T_4986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9568;
  reg [31:0] _T_4986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9569;
  reg [31:0] _T_4987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9570;
  reg [31:0] _T_4987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9571;
  reg [31:0] _T_4988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9572;
  reg [31:0] _T_4988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9573;
  reg [31:0] _T_4989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9574;
  reg [31:0] _T_4989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9575;
  reg [31:0] _T_4990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9576;
  reg [31:0] _T_4990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9577;
  reg [31:0] _T_4991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9578;
  reg [31:0] _T_4991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9579;
  reg [31:0] _T_4992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9580;
  reg [31:0] _T_4992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9581;
  reg [31:0] _T_4993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9582;
  reg [31:0] _T_4993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9583;
  reg [31:0] _T_4994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9584;
  reg [31:0] _T_4994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9585;
  reg [31:0] _T_4995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9586;
  reg [31:0] _T_4995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9587;
  reg [31:0] _T_4996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9588;
  reg [31:0] _T_4996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9589;
  reg [31:0] _T_4997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9590;
  reg [31:0] _T_4997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9591;
  reg [31:0] _T_4998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9592;
  reg [31:0] _T_4998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9593;
  reg [31:0] _T_4999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9594;
  reg [31:0] _T_4999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9595;
  reg [31:0] _T_5000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9596;
  reg [31:0] _T_5000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9597;
  reg [31:0] _T_5001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9598;
  reg [31:0] _T_5001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9599;
  reg [31:0] _T_5002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9600;
  reg [31:0] _T_5002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9601;
  reg [31:0] _T_5003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9602;
  reg [31:0] _T_5003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9603;
  reg [31:0] _T_5004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9604;
  reg [31:0] _T_5004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9605;
  reg [31:0] _T_5005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9606;
  reg [31:0] _T_5005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9607;
  reg [31:0] _T_5006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9608;
  reg [31:0] _T_5006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9609;
  reg [31:0] _T_5007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9610;
  reg [31:0] _T_5007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9611;
  reg [31:0] _T_5008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9612;
  reg [31:0] _T_5008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9613;
  reg [31:0] _T_5009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9614;
  reg [31:0] _T_5009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9615;
  reg [31:0] _T_5010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9616;
  reg [31:0] _T_5010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9617;
  reg [31:0] _T_5011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9618;
  reg [31:0] _T_5011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9619;
  reg [31:0] _T_5012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9620;
  reg [31:0] _T_5012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9621;
  reg [31:0] _T_5013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9622;
  reg [31:0] _T_5013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9623;
  reg [31:0] _T_5014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9624;
  reg [31:0] _T_5014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9625;
  reg [31:0] _T_5015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9626;
  reg [31:0] _T_5015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9627;
  reg [31:0] _T_5016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9628;
  reg [31:0] _T_5016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9629;
  reg [31:0] _T_5017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9630;
  reg [31:0] _T_5017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9631;
  reg [31:0] _T_5018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9632;
  reg [31:0] _T_5018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9633;
  reg [31:0] _T_5019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9634;
  reg [31:0] _T_5019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9635;
  reg [31:0] _T_5020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9636;
  reg [31:0] _T_5020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9637;
  reg [31:0] _T_5021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9638;
  reg [31:0] _T_5021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9639;
  reg [31:0] _T_5022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9640;
  reg [31:0] _T_5022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9641;
  reg [31:0] _T_5023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9642;
  reg [31:0] _T_5023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9643;
  reg [31:0] _T_5024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9644;
  reg [31:0] _T_5024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9645;
  reg [31:0] _T_5025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9646;
  reg [31:0] _T_5025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9647;
  reg [31:0] _T_5026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9648;
  reg [31:0] _T_5026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9649;
  reg [31:0] _T_5027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9650;
  reg [31:0] _T_5027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9651;
  reg [31:0] _T_5028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9652;
  reg [31:0] _T_5028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9653;
  reg [31:0] _T_5029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9654;
  reg [31:0] _T_5029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9655;
  reg [31:0] _T_5030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9656;
  reg [31:0] _T_5030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9657;
  reg [31:0] _T_5031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9658;
  reg [31:0] _T_5031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9659;
  reg [31:0] _T_5032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9660;
  reg [31:0] _T_5032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9661;
  reg [31:0] _T_5033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9662;
  reg [31:0] _T_5033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9663;
  reg [31:0] _T_5034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9664;
  reg [31:0] _T_5034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9665;
  reg [31:0] _T_5035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9666;
  reg [31:0] _T_5035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9667;
  reg [31:0] _T_5036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9668;
  reg [31:0] _T_5036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9669;
  reg [31:0] _T_5037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9670;
  reg [31:0] _T_5037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9671;
  reg [31:0] _T_5038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9672;
  reg [31:0] _T_5038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9673;
  reg [31:0] _T_5039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9674;
  reg [31:0] _T_5039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9675;
  reg [31:0] _T_5040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9676;
  reg [31:0] _T_5040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9677;
  reg [31:0] _T_5041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9678;
  reg [31:0] _T_5041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9679;
  reg [31:0] _T_5042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9680;
  reg [31:0] _T_5042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9681;
  reg [31:0] _T_5043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9682;
  reg [31:0] _T_5043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9683;
  reg [31:0] _T_5044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9684;
  reg [31:0] _T_5044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9685;
  reg [31:0] _T_5045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9686;
  reg [31:0] _T_5045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9687;
  reg [31:0] _T_5046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9688;
  reg [31:0] _T_5046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9689;
  reg [31:0] _T_5047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9690;
  reg [31:0] _T_5047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9691;
  reg [31:0] _T_5048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9692;
  reg [31:0] _T_5048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9693;
  reg [31:0] _T_5049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9694;
  reg [31:0] _T_5049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9695;
  reg [31:0] _T_5050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9696;
  reg [31:0] _T_5050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9697;
  reg [31:0] _T_5051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9698;
  reg [31:0] _T_5051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9699;
  reg [31:0] _T_5052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9700;
  reg [31:0] _T_5052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9701;
  reg [31:0] _T_5053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9702;
  reg [31:0] _T_5053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9703;
  reg [31:0] _T_5054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9704;
  reg [31:0] _T_5054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9705;
  reg [31:0] _T_5055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9706;
  reg [31:0] _T_5055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9707;
  reg [31:0] _T_5056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9708;
  reg [31:0] _T_5056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9709;
  reg [31:0] _T_5057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9710;
  reg [31:0] _T_5057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9711;
  reg [31:0] _T_5058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9712;
  reg [31:0] _T_5058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9713;
  reg [31:0] _T_5059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9714;
  reg [31:0] _T_5059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9715;
  reg [31:0] _T_5060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9716;
  reg [31:0] _T_5060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9717;
  reg [31:0] _T_5061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9718;
  reg [31:0] _T_5061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9719;
  reg [31:0] _T_5062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9720;
  reg [31:0] _T_5062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9721;
  reg [31:0] _T_5063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9722;
  reg [31:0] _T_5063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9723;
  reg [31:0] _T_5064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9724;
  reg [31:0] _T_5064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9725;
  reg [31:0] _T_5065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9726;
  reg [31:0] _T_5065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9727;
  reg [31:0] _T_5066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9728;
  reg [31:0] _T_5066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9729;
  reg [31:0] _T_5067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9730;
  reg [31:0] _T_5067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9731;
  reg [31:0] _T_5068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9732;
  reg [31:0] _T_5068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9733;
  reg [31:0] _T_5069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9734;
  reg [31:0] _T_5069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9735;
  reg [31:0] _T_5070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9736;
  reg [31:0] _T_5070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9737;
  reg [31:0] _T_5071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9738;
  reg [31:0] _T_5071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9739;
  reg [31:0] _T_5072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9740;
  reg [31:0] _T_5072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9741;
  reg [31:0] _T_5073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9742;
  reg [31:0] _T_5073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9743;
  reg [31:0] _T_5074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9744;
  reg [31:0] _T_5074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9745;
  reg [31:0] _T_5075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9746;
  reg [31:0] _T_5075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9747;
  reg [31:0] _T_5076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9748;
  reg [31:0] _T_5076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9749;
  reg [31:0] _T_5077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9750;
  reg [31:0] _T_5077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9751;
  reg [31:0] _T_5078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9752;
  reg [31:0] _T_5078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9753;
  reg [31:0] _T_5079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9754;
  reg [31:0] _T_5079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9755;
  reg [31:0] _T_5080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9756;
  reg [31:0] _T_5080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9757;
  reg [31:0] _T_5081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9758;
  reg [31:0] _T_5081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9759;
  reg [31:0] _T_5082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9760;
  reg [31:0] _T_5082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9761;
  reg [31:0] _T_5083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9762;
  reg [31:0] _T_5083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9763;
  reg [31:0] _T_5084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9764;
  reg [31:0] _T_5084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9765;
  reg [31:0] _T_5085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9766;
  reg [31:0] _T_5085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9767;
  reg [31:0] _T_5086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9768;
  reg [31:0] _T_5086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9769;
  reg [31:0] _T_5087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9770;
  reg [31:0] _T_5087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9771;
  reg [31:0] _T_5088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9772;
  reg [31:0] _T_5088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9773;
  reg [31:0] _T_5089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9774;
  reg [31:0] _T_5089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9775;
  reg [31:0] _T_5090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9776;
  reg [31:0] _T_5090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9777;
  reg [31:0] _T_5091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9778;
  reg [31:0] _T_5091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9779;
  reg [31:0] _T_5092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9780;
  reg [31:0] _T_5092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9781;
  reg [31:0] _T_5093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9782;
  reg [31:0] _T_5093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9783;
  reg [31:0] _T_5094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9784;
  reg [31:0] _T_5094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9785;
  reg [31:0] _T_5095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9786;
  reg [31:0] _T_5095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9787;
  reg [31:0] _T_5096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9788;
  reg [31:0] _T_5096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9789;
  reg [31:0] _T_5097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9790;
  reg [31:0] _T_5097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9791;
  reg [31:0] _T_5098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9792;
  reg [31:0] _T_5098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9793;
  reg [31:0] _T_5099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9794;
  reg [31:0] _T_5099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9795;
  reg [31:0] _T_5100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9796;
  reg [31:0] _T_5100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9797;
  reg [31:0] _T_5101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9798;
  reg [31:0] _T_5101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9799;
  reg [31:0] _T_5102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9800;
  reg [31:0] _T_5102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9801;
  reg [31:0] _T_5103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9802;
  reg [31:0] _T_5103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9803;
  reg [31:0] _T_5104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9804;
  reg [31:0] _T_5104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9805;
  reg [31:0] _T_5105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9806;
  reg [31:0] _T_5105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9807;
  reg [31:0] _T_5106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9808;
  reg [31:0] _T_5106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9809;
  reg [31:0] _T_5107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9810;
  reg [31:0] _T_5107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9811;
  reg [31:0] _T_5108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9812;
  reg [31:0] _T_5108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9813;
  reg [31:0] _T_5109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9814;
  reg [31:0] _T_5109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9815;
  reg [31:0] _T_5110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9816;
  reg [31:0] _T_5110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9817;
  reg [31:0] _T_5111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9818;
  reg [31:0] _T_5111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9819;
  reg [31:0] _T_5112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9820;
  reg [31:0] _T_5112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9821;
  reg [31:0] _T_5113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9822;
  reg [31:0] _T_5113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9823;
  reg [31:0] _T_5114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9824;
  reg [31:0] _T_5114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9825;
  reg [31:0] _T_5115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9826;
  reg [31:0] _T_5115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9827;
  reg [31:0] _T_5116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9828;
  reg [31:0] _T_5116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9829;
  reg [31:0] _T_5117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9830;
  reg [31:0] _T_5117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9831;
  reg [31:0] _T_5118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9832;
  reg [31:0] _T_5118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9833;
  reg [31:0] _T_5119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9834;
  reg [31:0] _T_5119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9835;
  reg [31:0] _T_5120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9836;
  reg [31:0] _T_5120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9837;
  reg [31:0] _T_5121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9838;
  reg [31:0] _T_5121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9839;
  reg [31:0] _T_5122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9840;
  reg [31:0] _T_5122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9841;
  reg [31:0] _T_5123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9842;
  reg [31:0] _T_5123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9843;
  reg [31:0] _T_5124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9844;
  reg [31:0] _T_5124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9845;
  reg [31:0] _T_5125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9846;
  reg [31:0] _T_5125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9847;
  reg [31:0] _T_5126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9848;
  reg [31:0] _T_5126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9849;
  reg [31:0] _T_5127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9850;
  reg [31:0] _T_5127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9851;
  reg [31:0] _T_5128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9852;
  reg [31:0] _T_5128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9853;
  reg [31:0] _T_5129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9854;
  reg [31:0] _T_5129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9855;
  reg [31:0] _T_5130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9856;
  reg [31:0] _T_5130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9857;
  reg [31:0] _T_5131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9858;
  reg [31:0] _T_5131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9859;
  reg [31:0] _T_5132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9860;
  reg [31:0] _T_5132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9861;
  reg [31:0] _T_5133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9862;
  reg [31:0] _T_5133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9863;
  reg [31:0] _T_5134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9864;
  reg [31:0] _T_5134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9865;
  reg [31:0] _T_5135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9866;
  reg [31:0] _T_5135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9867;
  reg [31:0] _T_5136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9868;
  reg [31:0] _T_5136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9869;
  reg [31:0] _T_5137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9870;
  reg [31:0] _T_5137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9871;
  reg [31:0] _T_5138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9872;
  reg [31:0] _T_5138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9873;
  reg [31:0] _T_5139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9874;
  reg [31:0] _T_5139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9875;
  reg [31:0] _T_5140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9876;
  reg [31:0] _T_5140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9877;
  reg [31:0] _T_5141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9878;
  reg [31:0] _T_5141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9879;
  reg [31:0] _T_5142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9880;
  reg [31:0] _T_5142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9881;
  reg [31:0] _T_5143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9882;
  reg [31:0] _T_5143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9883;
  reg [31:0] _T_5144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9884;
  reg [31:0] _T_5144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9885;
  reg [31:0] _T_5145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9886;
  reg [31:0] _T_5145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9887;
  reg [31:0] _T_5146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9888;
  reg [31:0] _T_5146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9889;
  reg [31:0] _T_5147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9890;
  reg [31:0] _T_5147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9891;
  reg [31:0] _T_5148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9892;
  reg [31:0] _T_5148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9893;
  reg [31:0] _T_5149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9894;
  reg [31:0] _T_5149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9895;
  reg [31:0] _T_5150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9896;
  reg [31:0] _T_5150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9897;
  reg [31:0] _T_5151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9898;
  reg [31:0] _T_5151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9899;
  reg [31:0] _T_5152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9900;
  reg [31:0] _T_5152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9901;
  reg [31:0] _T_5153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9902;
  reg [31:0] _T_5153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9903;
  reg [31:0] _T_5154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9904;
  reg [31:0] _T_5154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9905;
  reg [31:0] _T_5155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9906;
  reg [31:0] _T_5155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9907;
  reg [31:0] _T_5156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9908;
  reg [31:0] _T_5156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9909;
  reg [31:0] _T_5157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9910;
  reg [31:0] _T_5157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9911;
  reg [31:0] _T_5158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9912;
  reg [31:0] _T_5158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9913;
  reg [31:0] _T_5159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9914;
  reg [31:0] _T_5159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9915;
  reg [31:0] _T_5160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9916;
  reg [31:0] _T_5160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9917;
  reg [31:0] _T_5161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9918;
  reg [31:0] _T_5161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9919;
  reg [31:0] _T_5162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9920;
  reg [31:0] _T_5162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9921;
  reg [31:0] _T_5163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9922;
  reg [31:0] _T_5163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9923;
  reg [31:0] _T_5164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9924;
  reg [31:0] _T_5164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9925;
  reg [31:0] _T_5165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9926;
  reg [31:0] _T_5165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9927;
  reg [31:0] _T_5166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9928;
  reg [31:0] _T_5166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9929;
  reg [31:0] _T_5167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9930;
  reg [31:0] _T_5167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9931;
  reg [31:0] _T_5168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9932;
  reg [31:0] _T_5168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9933;
  reg [31:0] _T_5169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9934;
  reg [31:0] _T_5169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9935;
  reg [31:0] _T_5170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9936;
  reg [31:0] _T_5170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9937;
  reg [31:0] _T_5171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9938;
  reg [31:0] _T_5171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9939;
  reg [31:0] _T_5172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9940;
  reg [31:0] _T_5172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9941;
  reg [31:0] _T_5173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9942;
  reg [31:0] _T_5173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9943;
  reg [31:0] _T_5174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9944;
  reg [31:0] _T_5174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9945;
  reg [31:0] _T_5175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9946;
  reg [31:0] _T_5175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9947;
  reg [31:0] _T_5176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9948;
  reg [31:0] _T_5176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9949;
  reg [31:0] _T_5177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9950;
  reg [31:0] _T_5177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9951;
  reg [31:0] _T_5178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9952;
  reg [31:0] _T_5178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9953;
  reg [31:0] _T_5179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9954;
  reg [31:0] _T_5179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9955;
  reg [31:0] _T_5180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9956;
  reg [31:0] _T_5180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9957;
  reg [31:0] _T_5181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9958;
  reg [31:0] _T_5181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9959;
  reg [31:0] _T_5182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9960;
  reg [31:0] _T_5182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9961;
  reg [31:0] _T_5183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9962;
  reg [31:0] _T_5183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9963;
  reg [31:0] _T_5184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9964;
  reg [31:0] _T_5184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9965;
  reg [31:0] _T_5185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9966;
  reg [31:0] _T_5185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9967;
  reg [31:0] _T_5186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9968;
  reg [31:0] _T_5186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9969;
  reg [31:0] _T_5187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9970;
  reg [31:0] _T_5187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9971;
  reg [31:0] _T_5188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9972;
  reg [31:0] _T_5188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9973;
  reg [31:0] _T_5189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9974;
  reg [31:0] _T_5189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9975;
  reg [31:0] _T_5190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9976;
  reg [31:0] _T_5190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9977;
  reg [31:0] _T_5191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9978;
  reg [31:0] _T_5191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9979;
  reg [31:0] _T_5192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9980;
  reg [31:0] _T_5192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9981;
  reg [31:0] _T_5193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9982;
  reg [31:0] _T_5193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9983;
  reg [31:0] _T_5194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9984;
  reg [31:0] _T_5194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9985;
  reg [31:0] _T_5195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9986;
  reg [31:0] _T_5195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9987;
  reg [31:0] _T_5196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9988;
  reg [31:0] _T_5196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9989;
  reg [31:0] _T_5197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9990;
  reg [31:0] _T_5197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9991;
  reg [31:0] _T_5198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9992;
  reg [31:0] _T_5198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9993;
  reg [31:0] _T_5199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9994;
  reg [31:0] _T_5199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9995;
  reg [31:0] _T_5200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9996;
  reg [31:0] _T_5200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9997;
  reg [31:0] _T_5201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9998;
  reg [31:0] _T_5201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9999;
  reg [31:0] _T_5202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10000;
  reg [31:0] _T_5202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10001;
  reg [31:0] _T_5203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10002;
  reg [31:0] _T_5203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10003;
  reg [31:0] _T_5204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10004;
  reg [31:0] _T_5204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10005;
  reg [31:0] _T_5205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10006;
  reg [31:0] _T_5205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10007;
  reg [31:0] _T_5206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10008;
  reg [31:0] _T_5206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10009;
  reg [31:0] _T_5207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10010;
  reg [31:0] _T_5207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10011;
  reg [31:0] _T_5208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10012;
  reg [31:0] _T_5208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10013;
  reg [31:0] _T_5209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10014;
  reg [31:0] _T_5209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10015;
  reg [31:0] _T_5210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10016;
  reg [31:0] _T_5210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10017;
  reg [31:0] _T_5211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10018;
  reg [31:0] _T_5211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10019;
  reg [31:0] _T_5212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10020;
  reg [31:0] _T_5212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10021;
  reg [31:0] _T_5213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10022;
  reg [31:0] _T_5213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10023;
  reg [31:0] _T_5214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10024;
  reg [31:0] _T_5214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10025;
  reg [31:0] _T_5215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10026;
  reg [31:0] _T_5215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10027;
  reg [31:0] _T_5216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10028;
  reg [31:0] _T_5216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10029;
  reg [31:0] _T_5217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10030;
  reg [31:0] _T_5217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10031;
  reg [31:0] _T_5218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10032;
  reg [31:0] _T_5218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10033;
  reg [31:0] _T_5219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10034;
  reg [31:0] _T_5219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10035;
  reg [31:0] _T_5220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10036;
  reg [31:0] _T_5220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10037;
  reg [31:0] _T_5221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10038;
  reg [31:0] _T_5221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10039;
  reg [31:0] _T_5222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10040;
  reg [31:0] _T_5222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10041;
  reg [31:0] _T_5223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10042;
  reg [31:0] _T_5223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10043;
  reg [31:0] _T_5224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10044;
  reg [31:0] _T_5224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10045;
  reg [31:0] _T_5225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10046;
  reg [31:0] _T_5225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10047;
  reg [31:0] _T_5226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10048;
  reg [31:0] _T_5226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10049;
  reg [31:0] _T_5227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10050;
  reg [31:0] _T_5227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10051;
  reg [31:0] _T_5228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10052;
  reg [31:0] _T_5228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10053;
  reg [31:0] _T_5229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10054;
  reg [31:0] _T_5229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10055;
  reg [31:0] _T_5230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10056;
  reg [31:0] _T_5230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10057;
  reg [31:0] _T_5231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10058;
  reg [31:0] _T_5231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10059;
  reg [31:0] _T_5232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10060;
  reg [31:0] _T_5232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10061;
  reg [31:0] _T_5233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10062;
  reg [31:0] _T_5233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10063;
  reg [31:0] _T_5234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10064;
  reg [31:0] _T_5234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10065;
  reg [31:0] _T_5235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10066;
  reg [31:0] _T_5235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10067;
  reg [31:0] _T_5236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10068;
  reg [31:0] _T_5236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10069;
  reg [31:0] _T_5237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10070;
  reg [31:0] _T_5237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10071;
  reg [31:0] _T_5238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10072;
  reg [31:0] _T_5238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10073;
  reg [31:0] _T_5239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10074;
  reg [31:0] _T_5239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10075;
  reg [31:0] _T_5240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10076;
  reg [31:0] _T_5240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10077;
  reg [31:0] _T_5241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10078;
  reg [31:0] _T_5241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10079;
  reg [31:0] _T_5242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10080;
  reg [31:0] _T_5242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10081;
  reg [31:0] _T_5243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10082;
  reg [31:0] _T_5243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10083;
  reg [31:0] _T_5244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10084;
  reg [31:0] _T_5244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10085;
  reg [31:0] _T_5245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10086;
  reg [31:0] _T_5245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10087;
  reg [31:0] _T_5246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10088;
  reg [31:0] _T_5246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10089;
  reg [31:0] _T_5247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10090;
  reg [31:0] _T_5247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10091;
  reg [31:0] _T_5248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10092;
  reg [31:0] _T_5248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10093;
  reg [31:0] _T_5249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10094;
  reg [31:0] _T_5249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10095;
  reg [31:0] _T_5250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10096;
  reg [31:0] _T_5250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10097;
  reg [31:0] _T_5251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10098;
  reg [31:0] _T_5251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10099;
  reg [31:0] _T_5252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10100;
  reg [31:0] _T_5252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10101;
  reg [31:0] _T_5253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10102;
  reg [31:0] _T_5253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10103;
  reg [31:0] _T_5254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10104;
  reg [31:0] _T_5254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10105;
  reg [31:0] _T_5255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10106;
  reg [31:0] _T_5255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10107;
  reg [31:0] _T_5256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10108;
  reg [31:0] _T_5256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10109;
  reg [31:0] _T_5257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10110;
  reg [31:0] _T_5257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10111;
  reg [31:0] _T_5258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10112;
  reg [31:0] _T_5258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10113;
  reg [31:0] _T_5259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10114;
  reg [31:0] _T_5259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10115;
  reg [31:0] _T_5260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10116;
  reg [31:0] _T_5260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10117;
  reg [31:0] _T_5261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10118;
  reg [31:0] _T_5261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10119;
  reg [31:0] _T_5262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10120;
  reg [31:0] _T_5262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10121;
  reg [31:0] _T_5263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10122;
  reg [31:0] _T_5263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10123;
  reg [31:0] _T_5264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10124;
  reg [31:0] _T_5264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10125;
  reg [31:0] _T_5265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10126;
  reg [31:0] _T_5265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10127;
  reg [31:0] _T_5266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10128;
  reg [31:0] _T_5266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10129;
  reg [31:0] _T_5267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10130;
  reg [31:0] _T_5267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10131;
  reg [31:0] _T_5268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10132;
  reg [31:0] _T_5268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10133;
  reg [31:0] _T_5269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10134;
  reg [31:0] _T_5269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10135;
  reg [31:0] _T_5270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10136;
  reg [31:0] _T_5270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10137;
  reg [31:0] _T_5271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10138;
  reg [31:0] _T_5271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10139;
  reg [31:0] _T_5272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10140;
  reg [31:0] _T_5272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10141;
  reg [31:0] _T_5273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10142;
  reg [31:0] _T_5273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10143;
  reg [31:0] _T_5274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10144;
  reg [31:0] _T_5274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10145;
  reg [31:0] _T_5275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10146;
  reg [31:0] _T_5275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10147;
  reg [31:0] _T_5276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10148;
  reg [31:0] _T_5276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10149;
  reg [31:0] _T_5277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10150;
  reg [31:0] _T_5277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10151;
  reg [31:0] _T_5278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10152;
  reg [31:0] _T_5278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10153;
  reg [31:0] _T_5279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10154;
  reg [31:0] _T_5279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10155;
  reg [31:0] _T_5280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10156;
  reg [31:0] _T_5280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10157;
  reg [31:0] _T_5281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10158;
  reg [31:0] _T_5281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10159;
  reg [31:0] _T_5282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10160;
  reg [31:0] _T_5282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10161;
  reg [31:0] _T_5283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10162;
  reg [31:0] _T_5283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10163;
  reg [31:0] _T_5284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10164;
  reg [31:0] _T_5284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10165;
  reg [31:0] _T_5285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10166;
  reg [31:0] _T_5285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10167;
  reg [31:0] _T_5286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10168;
  reg [31:0] _T_5286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10169;
  reg [31:0] _T_5287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10170;
  reg [31:0] _T_5287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10171;
  reg [31:0] _T_5288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10172;
  reg [31:0] _T_5288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10173;
  reg [31:0] _T_5289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10174;
  reg [31:0] _T_5289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10175;
  reg [31:0] _T_5290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10176;
  reg [31:0] _T_5290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10177;
  reg [31:0] _T_5291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10178;
  reg [31:0] _T_5291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10179;
  reg [31:0] _T_5292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10180;
  reg [31:0] _T_5292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10181;
  reg [31:0] _T_5293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10182;
  reg [31:0] _T_5293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10183;
  reg [31:0] _T_5294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10184;
  reg [31:0] _T_5294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10185;
  reg [31:0] _T_5295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10186;
  reg [31:0] _T_5295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10187;
  reg [31:0] _T_5296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10188;
  reg [31:0] _T_5296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10189;
  reg [31:0] _T_5297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10190;
  reg [31:0] _T_5297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10191;
  reg [31:0] _T_5298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10192;
  reg [31:0] _T_5298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10193;
  reg [31:0] _T_5299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10194;
  reg [31:0] _T_5299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10195;
  reg [31:0] _T_5300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10196;
  reg [31:0] _T_5300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10197;
  reg [31:0] _T_5301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10198;
  reg [31:0] _T_5301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10199;
  reg [31:0] _T_5302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10200;
  reg [31:0] _T_5302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10201;
  reg [31:0] _T_5303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10202;
  reg [31:0] _T_5303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10203;
  reg [31:0] _T_5304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10204;
  reg [31:0] _T_5304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10205;
  reg [31:0] _T_5305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10206;
  reg [31:0] _T_5305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10207;
  reg [31:0] _T_5306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10208;
  reg [31:0] _T_5306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10209;
  reg [31:0] _T_5307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10210;
  reg [31:0] _T_5307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10211;
  reg [31:0] _T_5308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10212;
  reg [31:0] _T_5308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10213;
  reg [31:0] _T_5309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10214;
  reg [31:0] _T_5309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10215;
  reg [31:0] _T_5310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10216;
  reg [31:0] _T_5310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10217;
  reg [31:0] _T_5311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10218;
  reg [31:0] _T_5311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10219;
  reg [31:0] _T_5312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10220;
  reg [31:0] _T_5312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10221;
  reg [31:0] _T_5313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10222;
  reg [31:0] _T_5313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10223;
  reg [31:0] _T_5314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10224;
  reg [31:0] _T_5314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10225;
  reg [31:0] _T_5315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10226;
  reg [31:0] _T_5315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10227;
  reg [31:0] _T_5316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10228;
  reg [31:0] _T_5316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10229;
  reg [31:0] _T_5317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10230;
  reg [31:0] _T_5317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10231;
  reg [31:0] _T_5318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10232;
  reg [31:0] _T_5318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10233;
  reg [31:0] _T_5319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10234;
  reg [31:0] _T_5319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10235;
  reg [31:0] _T_5320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10236;
  reg [31:0] _T_5320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10237;
  reg [31:0] _T_5321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10238;
  reg [31:0] _T_5321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10239;
  reg [31:0] _T_5322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10240;
  reg [31:0] _T_5322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10241;
  reg [31:0] _T_5325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10242;
  reg [31:0] _T_5325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10243;
  reg [31:0] _T_5326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10244;
  reg [31:0] _T_5326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10245;
  reg [31:0] _T_5327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10246;
  reg [31:0] _T_5327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10247;
  reg [31:0] _T_5328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10248;
  reg [31:0] _T_5328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10249;
  reg [31:0] _T_5329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10250;
  reg [31:0] _T_5329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10251;
  reg [31:0] _T_5330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10252;
  reg [31:0] _T_5330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10253;
  reg [31:0] _T_5331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10254;
  reg [31:0] _T_5331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10255;
  reg [31:0] _T_5332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10256;
  reg [31:0] _T_5332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10257;
  reg [31:0] _T_5333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10258;
  reg [31:0] _T_5333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10259;
  reg [31:0] _T_5334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10260;
  reg [31:0] _T_5334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10261;
  reg [31:0] _T_5335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10262;
  reg [31:0] _T_5335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10263;
  reg [31:0] _T_5336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10264;
  reg [31:0] _T_5336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10265;
  reg [31:0] _T_5337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10266;
  reg [31:0] _T_5337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10267;
  reg [31:0] _T_5338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10268;
  reg [31:0] _T_5338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10269;
  reg [31:0] _T_5339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10270;
  reg [31:0] _T_5339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10271;
  reg [31:0] _T_5340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10272;
  reg [31:0] _T_5340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10273;
  reg [31:0] _T_5341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10274;
  reg [31:0] _T_5341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10275;
  reg [31:0] _T_5342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10276;
  reg [31:0] _T_5342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10277;
  reg [31:0] _T_5343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10278;
  reg [31:0] _T_5343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10279;
  reg [31:0] _T_5344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10280;
  reg [31:0] _T_5344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10281;
  reg [31:0] _T_5345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10282;
  reg [31:0] _T_5345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10283;
  reg [31:0] _T_5346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10284;
  reg [31:0] _T_5346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10285;
  reg [31:0] _T_5347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10286;
  reg [31:0] _T_5347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10287;
  reg [31:0] _T_5348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10288;
  reg [31:0] _T_5348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10289;
  reg [31:0] _T_5349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10290;
  reg [31:0] _T_5349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10291;
  reg [31:0] _T_5350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10292;
  reg [31:0] _T_5350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10293;
  reg [31:0] _T_5351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10294;
  reg [31:0] _T_5351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10295;
  reg [31:0] _T_5352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10296;
  reg [31:0] _T_5352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10297;
  reg [31:0] _T_5353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10298;
  reg [31:0] _T_5353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10299;
  reg [31:0] _T_5354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10300;
  reg [31:0] _T_5354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10301;
  reg [31:0] _T_5355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10302;
  reg [31:0] _T_5355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10303;
  reg [31:0] _T_5356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10304;
  reg [31:0] _T_5356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10305;
  reg [31:0] _T_5357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10306;
  reg [31:0] _T_5357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10307;
  reg [31:0] _T_5358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10308;
  reg [31:0] _T_5358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10309;
  reg [31:0] _T_5359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10310;
  reg [31:0] _T_5359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10311;
  reg [31:0] _T_5360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10312;
  reg [31:0] _T_5360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10313;
  reg [31:0] _T_5361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10314;
  reg [31:0] _T_5361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10315;
  reg [31:0] _T_5362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10316;
  reg [31:0] _T_5362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10317;
  reg [31:0] _T_5363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10318;
  reg [31:0] _T_5363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10319;
  reg [31:0] _T_5364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10320;
  reg [31:0] _T_5364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10321;
  reg [31:0] _T_5365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10322;
  reg [31:0] _T_5365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10323;
  reg [31:0] _T_5366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10324;
  reg [31:0] _T_5366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10325;
  reg [31:0] _T_5367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10326;
  reg [31:0] _T_5367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10327;
  reg [31:0] _T_5368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10328;
  reg [31:0] _T_5368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10329;
  reg [31:0] _T_5369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10330;
  reg [31:0] _T_5369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10331;
  reg [31:0] _T_5370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10332;
  reg [31:0] _T_5370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10333;
  reg [31:0] _T_5371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10334;
  reg [31:0] _T_5371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10335;
  reg [31:0] _T_5372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10336;
  reg [31:0] _T_5372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10337;
  reg [31:0] _T_5373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10338;
  reg [31:0] _T_5373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10339;
  reg [31:0] _T_5374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10340;
  reg [31:0] _T_5374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10341;
  reg [31:0] _T_5375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10342;
  reg [31:0] _T_5375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10343;
  reg [31:0] _T_5376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10344;
  reg [31:0] _T_5376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10345;
  reg [31:0] _T_5377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10346;
  reg [31:0] _T_5377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10347;
  reg [31:0] _T_5378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10348;
  reg [31:0] _T_5378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10349;
  reg [31:0] _T_5379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10350;
  reg [31:0] _T_5379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10351;
  reg [31:0] _T_5380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10352;
  reg [31:0] _T_5380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10353;
  reg [31:0] _T_5381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10354;
  reg [31:0] _T_5381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10355;
  reg [31:0] _T_5382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10356;
  reg [31:0] _T_5382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10357;
  reg [31:0] _T_5383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10358;
  reg [31:0] _T_5383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10359;
  reg [31:0] _T_5384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10360;
  reg [31:0] _T_5384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10361;
  reg [31:0] _T_5385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10362;
  reg [31:0] _T_5385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10363;
  reg [31:0] _T_5386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10364;
  reg [31:0] _T_5386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10365;
  reg [31:0] _T_5387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10366;
  reg [31:0] _T_5387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10367;
  reg [31:0] _T_5388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10368;
  reg [31:0] _T_5388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10369;
  reg [31:0] _T_5389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10370;
  reg [31:0] _T_5389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10371;
  reg [31:0] _T_5390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10372;
  reg [31:0] _T_5390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10373;
  reg [31:0] _T_5391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10374;
  reg [31:0] _T_5391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10375;
  reg [31:0] _T_5392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10376;
  reg [31:0] _T_5392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10377;
  reg [31:0] _T_5393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10378;
  reg [31:0] _T_5393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10379;
  reg [31:0] _T_5394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10380;
  reg [31:0] _T_5394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10381;
  reg [31:0] _T_5395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10382;
  reg [31:0] _T_5395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10383;
  reg [31:0] _T_5396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10384;
  reg [31:0] _T_5396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10385;
  reg [31:0] _T_5397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10386;
  reg [31:0] _T_5397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10387;
  reg [31:0] _T_5398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10388;
  reg [31:0] _T_5398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10389;
  reg [31:0] _T_5399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10390;
  reg [31:0] _T_5399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10391;
  reg [31:0] _T_5400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10392;
  reg [31:0] _T_5400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10393;
  reg [31:0] _T_5401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10394;
  reg [31:0] _T_5401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10395;
  reg [31:0] _T_5402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10396;
  reg [31:0] _T_5402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10397;
  reg [31:0] _T_5403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10398;
  reg [31:0] _T_5403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10399;
  reg [31:0] _T_5404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10400;
  reg [31:0] _T_5404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10401;
  reg [31:0] _T_5405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10402;
  reg [31:0] _T_5405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10403;
  reg [31:0] _T_5406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10404;
  reg [31:0] _T_5406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10405;
  reg [31:0] _T_5407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10406;
  reg [31:0] _T_5407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10407;
  reg [31:0] _T_5408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10408;
  reg [31:0] _T_5408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10409;
  reg [31:0] _T_5409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10410;
  reg [31:0] _T_5409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10411;
  reg [31:0] _T_5410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10412;
  reg [31:0] _T_5410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10413;
  reg [31:0] _T_5411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10414;
  reg [31:0] _T_5411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10415;
  reg [31:0] _T_5412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10416;
  reg [31:0] _T_5412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10417;
  reg [31:0] _T_5413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10418;
  reg [31:0] _T_5413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10419;
  reg [31:0] _T_5414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10420;
  reg [31:0] _T_5414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10421;
  reg [31:0] _T_5415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10422;
  reg [31:0] _T_5415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10423;
  reg [31:0] _T_5416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10424;
  reg [31:0] _T_5416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10425;
  reg [31:0] _T_5417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10426;
  reg [31:0] _T_5417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10427;
  reg [31:0] _T_5418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10428;
  reg [31:0] _T_5418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10429;
  reg [31:0] _T_5419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10430;
  reg [31:0] _T_5419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10431;
  reg [31:0] _T_5420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10432;
  reg [31:0] _T_5420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10433;
  reg [31:0] _T_5421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10434;
  reg [31:0] _T_5421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10435;
  reg [31:0] _T_5422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10436;
  reg [31:0] _T_5422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10437;
  reg [31:0] _T_5423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10438;
  reg [31:0] _T_5423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10439;
  reg [31:0] _T_5424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10440;
  reg [31:0] _T_5424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10441;
  reg [31:0] _T_5425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10442;
  reg [31:0] _T_5425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10443;
  reg [31:0] _T_5426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10444;
  reg [31:0] _T_5426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10445;
  reg [31:0] _T_5427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10446;
  reg [31:0] _T_5427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10447;
  reg [31:0] _T_5428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10448;
  reg [31:0] _T_5428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10449;
  reg [31:0] _T_5429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10450;
  reg [31:0] _T_5429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10451;
  reg [31:0] _T_5430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10452;
  reg [31:0] _T_5430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10453;
  reg [31:0] _T_5431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10454;
  reg [31:0] _T_5431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10455;
  reg [31:0] _T_5432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10456;
  reg [31:0] _T_5432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10457;
  reg [31:0] _T_5433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10458;
  reg [31:0] _T_5433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10459;
  reg [31:0] _T_5434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10460;
  reg [31:0] _T_5434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10461;
  reg [31:0] _T_5435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10462;
  reg [31:0] _T_5435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10463;
  reg [31:0] _T_5436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10464;
  reg [31:0] _T_5436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10465;
  reg [31:0] _T_5437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10466;
  reg [31:0] _T_5437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10467;
  reg [31:0] _T_5438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10468;
  reg [31:0] _T_5438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10469;
  reg [31:0] _T_5439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10470;
  reg [31:0] _T_5439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10471;
  reg [31:0] _T_5440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10472;
  reg [31:0] _T_5440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10473;
  reg [31:0] _T_5441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10474;
  reg [31:0] _T_5441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10475;
  reg [31:0] _T_5442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10476;
  reg [31:0] _T_5442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10477;
  reg [31:0] _T_5443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10478;
  reg [31:0] _T_5443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10479;
  reg [31:0] _T_5444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10480;
  reg [31:0] _T_5444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10481;
  reg [31:0] _T_5445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10482;
  reg [31:0] _T_5445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10483;
  reg [31:0] _T_5446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10484;
  reg [31:0] _T_5446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10485;
  reg [31:0] _T_5447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10486;
  reg [31:0] _T_5447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10487;
  reg [31:0] _T_5448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10488;
  reg [31:0] _T_5448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10489;
  reg [31:0] _T_5449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10490;
  reg [31:0] _T_5449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10491;
  reg [31:0] _T_5450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10492;
  reg [31:0] _T_5450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10493;
  reg [31:0] _T_5451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10494;
  reg [31:0] _T_5451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10495;
  reg [31:0] _T_5452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10496;
  reg [31:0] _T_5452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10497;
  reg [31:0] _T_5453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10498;
  reg [31:0] _T_5453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10499;
  reg [31:0] _T_5454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10500;
  reg [31:0] _T_5454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10501;
  reg [31:0] _T_5455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10502;
  reg [31:0] _T_5455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10503;
  reg [31:0] _T_5456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10504;
  reg [31:0] _T_5456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10505;
  reg [31:0] _T_5457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10506;
  reg [31:0] _T_5457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10507;
  reg [31:0] _T_5458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10508;
  reg [31:0] _T_5458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10509;
  reg [31:0] _T_5459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10510;
  reg [31:0] _T_5459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10511;
  reg [31:0] _T_5460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10512;
  reg [31:0] _T_5460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10513;
  reg [31:0] _T_5461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10514;
  reg [31:0] _T_5461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10515;
  reg [31:0] _T_5462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10516;
  reg [31:0] _T_5462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10517;
  reg [31:0] _T_5463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10518;
  reg [31:0] _T_5463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10519;
  reg [31:0] _T_5464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10520;
  reg [31:0] _T_5464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10521;
  reg [31:0] _T_5465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10522;
  reg [31:0] _T_5465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10523;
  reg [31:0] _T_5466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10524;
  reg [31:0] _T_5466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10525;
  reg [31:0] _T_5467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10526;
  reg [31:0] _T_5467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10527;
  reg [31:0] _T_5468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10528;
  reg [31:0] _T_5468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10529;
  reg [31:0] _T_5469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10530;
  reg [31:0] _T_5469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10531;
  reg [31:0] _T_5470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10532;
  reg [31:0] _T_5470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10533;
  reg [31:0] _T_5471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10534;
  reg [31:0] _T_5471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10535;
  reg [31:0] _T_5472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10536;
  reg [31:0] _T_5472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10537;
  reg [31:0] _T_5473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10538;
  reg [31:0] _T_5473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10539;
  reg [31:0] _T_5474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10540;
  reg [31:0] _T_5474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10541;
  reg [31:0] _T_5475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10542;
  reg [31:0] _T_5475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10543;
  reg [31:0] _T_5476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10544;
  reg [31:0] _T_5476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10545;
  reg [31:0] _T_5477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10546;
  reg [31:0] _T_5477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10547;
  reg [31:0] _T_5478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10548;
  reg [31:0] _T_5478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10549;
  reg [31:0] _T_5479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10550;
  reg [31:0] _T_5479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10551;
  reg [31:0] _T_5480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10552;
  reg [31:0] _T_5480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10553;
  reg [31:0] _T_5481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10554;
  reg [31:0] _T_5481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10555;
  reg [31:0] _T_5482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10556;
  reg [31:0] _T_5482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10557;
  reg [31:0] _T_5483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10558;
  reg [31:0] _T_5483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10559;
  reg [31:0] _T_5484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10560;
  reg [31:0] _T_5484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10561;
  reg [31:0] _T_5485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10562;
  reg [31:0] _T_5485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10563;
  reg [31:0] _T_5486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10564;
  reg [31:0] _T_5486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10565;
  reg [31:0] _T_5487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10566;
  reg [31:0] _T_5487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10567;
  reg [31:0] _T_5488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10568;
  reg [31:0] _T_5488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10569;
  reg [31:0] _T_5489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10570;
  reg [31:0] _T_5489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10571;
  reg [31:0] _T_5490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10572;
  reg [31:0] _T_5490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10573;
  reg [31:0] _T_5491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10574;
  reg [31:0] _T_5491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10575;
  reg [31:0] _T_5492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10576;
  reg [31:0] _T_5492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10577;
  reg [31:0] _T_5493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10578;
  reg [31:0] _T_5493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10579;
  reg [31:0] _T_5494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10580;
  reg [31:0] _T_5494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10581;
  reg [31:0] _T_5495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10582;
  reg [31:0] _T_5495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10583;
  reg [31:0] _T_5496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10584;
  reg [31:0] _T_5496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10585;
  reg [31:0] _T_5497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10586;
  reg [31:0] _T_5497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10587;
  reg [31:0] _T_5498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10588;
  reg [31:0] _T_5498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10589;
  reg [31:0] _T_5499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10590;
  reg [31:0] _T_5499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10591;
  reg [31:0] _T_5500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10592;
  reg [31:0] _T_5500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10593;
  reg [31:0] _T_5501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10594;
  reg [31:0] _T_5501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10595;
  reg [31:0] _T_5502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10596;
  reg [31:0] _T_5502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10597;
  reg [31:0] _T_5503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10598;
  reg [31:0] _T_5503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10599;
  reg [31:0] _T_5504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10600;
  reg [31:0] _T_5504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10601;
  reg [31:0] _T_5505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10602;
  reg [31:0] _T_5505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10603;
  reg [31:0] _T_5506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10604;
  reg [31:0] _T_5506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10605;
  reg [31:0] _T_5507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10606;
  reg [31:0] _T_5507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10607;
  reg [31:0] _T_5508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10608;
  reg [31:0] _T_5508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10609;
  reg [31:0] _T_5509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10610;
  reg [31:0] _T_5509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10611;
  reg [31:0] _T_5510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10612;
  reg [31:0] _T_5510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10613;
  reg [31:0] _T_5511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10614;
  reg [31:0] _T_5511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10615;
  reg [31:0] _T_5512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10616;
  reg [31:0] _T_5512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10617;
  reg [31:0] _T_5513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10618;
  reg [31:0] _T_5513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10619;
  reg [31:0] _T_5514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10620;
  reg [31:0] _T_5514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10621;
  reg [31:0] _T_5515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10622;
  reg [31:0] _T_5515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10623;
  reg [31:0] _T_5516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10624;
  reg [31:0] _T_5516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10625;
  reg [31:0] _T_5517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10626;
  reg [31:0] _T_5517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10627;
  reg [31:0] _T_5518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10628;
  reg [31:0] _T_5518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10629;
  reg [31:0] _T_5519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10630;
  reg [31:0] _T_5519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10631;
  reg [31:0] _T_5520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10632;
  reg [31:0] _T_5520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10633;
  reg [31:0] _T_5521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10634;
  reg [31:0] _T_5521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10635;
  reg [31:0] _T_5522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10636;
  reg [31:0] _T_5522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10637;
  reg [31:0] _T_5523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10638;
  reg [31:0] _T_5523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10639;
  reg [31:0] _T_5524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10640;
  reg [31:0] _T_5524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10641;
  reg [31:0] _T_5525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10642;
  reg [31:0] _T_5525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10643;
  reg [31:0] _T_5526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10644;
  reg [31:0] _T_5526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10645;
  reg [31:0] _T_5527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10646;
  reg [31:0] _T_5527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10647;
  reg [31:0] _T_5528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10648;
  reg [31:0] _T_5528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10649;
  reg [31:0] _T_5529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10650;
  reg [31:0] _T_5529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10651;
  reg [31:0] _T_5530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10652;
  reg [31:0] _T_5530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10653;
  reg [31:0] _T_5531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10654;
  reg [31:0] _T_5531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10655;
  reg [31:0] _T_5532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10656;
  reg [31:0] _T_5532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10657;
  reg [31:0] _T_5533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10658;
  reg [31:0] _T_5533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10659;
  reg [31:0] _T_5534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10660;
  reg [31:0] _T_5534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10661;
  reg [31:0] _T_5535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10662;
  reg [31:0] _T_5535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10663;
  reg [31:0] _T_5536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10664;
  reg [31:0] _T_5536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10665;
  reg [31:0] _T_5537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10666;
  reg [31:0] _T_5537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10667;
  reg [31:0] _T_5538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10668;
  reg [31:0] _T_5538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10669;
  reg [31:0] _T_5539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10670;
  reg [31:0] _T_5539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10671;
  reg [31:0] _T_5540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10672;
  reg [31:0] _T_5540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10673;
  reg [31:0] _T_5541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10674;
  reg [31:0] _T_5541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10675;
  reg [31:0] _T_5542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10676;
  reg [31:0] _T_5542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10677;
  reg [31:0] _T_5543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10678;
  reg [31:0] _T_5543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10679;
  reg [31:0] _T_5544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10680;
  reg [31:0] _T_5544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10681;
  reg [31:0] _T_5545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10682;
  reg [31:0] _T_5545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10683;
  reg [31:0] _T_5546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10684;
  reg [31:0] _T_5546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10685;
  reg [31:0] _T_5547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10686;
  reg [31:0] _T_5547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10687;
  reg [31:0] _T_5548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10688;
  reg [31:0] _T_5548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10689;
  reg [31:0] _T_5549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10690;
  reg [31:0] _T_5549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10691;
  reg [31:0] _T_5550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10692;
  reg [31:0] _T_5550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10693;
  reg [31:0] _T_5551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10694;
  reg [31:0] _T_5551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10695;
  reg [31:0] _T_5552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10696;
  reg [31:0] _T_5552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10697;
  reg [31:0] _T_5553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10698;
  reg [31:0] _T_5553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10699;
  reg [31:0] _T_5554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10700;
  reg [31:0] _T_5554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10701;
  reg [31:0] _T_5555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10702;
  reg [31:0] _T_5555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10703;
  reg [31:0] _T_5556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10704;
  reg [31:0] _T_5556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10705;
  reg [31:0] _T_5557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10706;
  reg [31:0] _T_5557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10707;
  reg [31:0] _T_5558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10708;
  reg [31:0] _T_5558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10709;
  reg [31:0] _T_5559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10710;
  reg [31:0] _T_5559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10711;
  reg [31:0] _T_5560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10712;
  reg [31:0] _T_5560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10713;
  reg [31:0] _T_5561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10714;
  reg [31:0] _T_5561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10715;
  reg [31:0] _T_5562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10716;
  reg [31:0] _T_5562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10717;
  reg [31:0] _T_5563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10718;
  reg [31:0] _T_5563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10719;
  reg [31:0] _T_5564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10720;
  reg [31:0] _T_5564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10721;
  reg [31:0] _T_5565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10722;
  reg [31:0] _T_5565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10723;
  reg [31:0] _T_5566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10724;
  reg [31:0] _T_5566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10725;
  reg [31:0] _T_5567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10726;
  reg [31:0] _T_5567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10727;
  reg [31:0] _T_5568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10728;
  reg [31:0] _T_5568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10729;
  reg [31:0] _T_5569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10730;
  reg [31:0] _T_5569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10731;
  reg [31:0] _T_5570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10732;
  reg [31:0] _T_5570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10733;
  reg [31:0] _T_5571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10734;
  reg [31:0] _T_5571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10735;
  reg [31:0] _T_5572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10736;
  reg [31:0] _T_5572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10737;
  reg [31:0] _T_5573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10738;
  reg [31:0] _T_5573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10739;
  reg [31:0] _T_5574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10740;
  reg [31:0] _T_5574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10741;
  reg [31:0] _T_5575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10742;
  reg [31:0] _T_5575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10743;
  reg [31:0] _T_5576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10744;
  reg [31:0] _T_5576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10745;
  reg [31:0] _T_5577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10746;
  reg [31:0] _T_5577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10747;
  reg [31:0] _T_5578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10748;
  reg [31:0] _T_5578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10749;
  reg [31:0] _T_5579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10750;
  reg [31:0] _T_5579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10751;
  reg [31:0] _T_5580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10752;
  reg [31:0] _T_5580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10753;
  wire [31:0] _GEN_17922 = 8'h1 == cnt[7:0] ? $signed(32'shfffb) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17923 = 8'h2 == cnt[7:0] ? $signed(32'shffec) : $signed(_GEN_17922); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17924 = 8'h3 == cnt[7:0] ? $signed(32'shffd4) : $signed(_GEN_17923); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17925 = 8'h4 == cnt[7:0] ? $signed(32'shffb1) : $signed(_GEN_17924); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17926 = 8'h5 == cnt[7:0] ? $signed(32'shff85) : $signed(_GEN_17925); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17927 = 8'h6 == cnt[7:0] ? $signed(32'shff4e) : $signed(_GEN_17926); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17928 = 8'h7 == cnt[7:0] ? $signed(32'shff0e) : $signed(_GEN_17927); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17929 = 8'h8 == cnt[7:0] ? $signed(32'shfec4) : $signed(_GEN_17928); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17930 = 8'h9 == cnt[7:0] ? $signed(32'shfe71) : $signed(_GEN_17929); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17931 = 8'ha == cnt[7:0] ? $signed(32'shfe13) : $signed(_GEN_17930); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17932 = 8'hb == cnt[7:0] ? $signed(32'shfdac) : $signed(_GEN_17931); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17933 = 8'hc == cnt[7:0] ? $signed(32'shfd3b) : $signed(_GEN_17932); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17934 = 8'hd == cnt[7:0] ? $signed(32'shfcc0) : $signed(_GEN_17933); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17935 = 8'he == cnt[7:0] ? $signed(32'shfc3b) : $signed(_GEN_17934); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17936 = 8'hf == cnt[7:0] ? $signed(32'shfbad) : $signed(_GEN_17935); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17937 = 8'h10 == cnt[7:0] ? $signed(32'shfb15) : $signed(_GEN_17936); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17938 = 8'h11 == cnt[7:0] ? $signed(32'shfa73) : $signed(_GEN_17937); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17939 = 8'h12 == cnt[7:0] ? $signed(32'shf9c8) : $signed(_GEN_17938); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17940 = 8'h13 == cnt[7:0] ? $signed(32'shf913) : $signed(_GEN_17939); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17941 = 8'h14 == cnt[7:0] ? $signed(32'shf854) : $signed(_GEN_17940); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17942 = 8'h15 == cnt[7:0] ? $signed(32'shf78c) : $signed(_GEN_17941); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17943 = 8'h16 == cnt[7:0] ? $signed(32'shf6ba) : $signed(_GEN_17942); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17944 = 8'h17 == cnt[7:0] ? $signed(32'shf5df) : $signed(_GEN_17943); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17945 = 8'h18 == cnt[7:0] ? $signed(32'shf4fa) : $signed(_GEN_17944); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17946 = 8'h19 == cnt[7:0] ? $signed(32'shf40c) : $signed(_GEN_17945); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17947 = 8'h1a == cnt[7:0] ? $signed(32'shf314) : $signed(_GEN_17946); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17948 = 8'h1b == cnt[7:0] ? $signed(32'shf213) : $signed(_GEN_17947); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17949 = 8'h1c == cnt[7:0] ? $signed(32'shf109) : $signed(_GEN_17948); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17950 = 8'h1d == cnt[7:0] ? $signed(32'sheff5) : $signed(_GEN_17949); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17951 = 8'h1e == cnt[7:0] ? $signed(32'sheed9) : $signed(_GEN_17950); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17952 = 8'h1f == cnt[7:0] ? $signed(32'shedb3) : $signed(_GEN_17951); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17953 = 8'h20 == cnt[7:0] ? $signed(32'shec83) : $signed(_GEN_17952); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17954 = 8'h21 == cnt[7:0] ? $signed(32'sheb4b) : $signed(_GEN_17953); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17955 = 8'h22 == cnt[7:0] ? $signed(32'shea0a) : $signed(_GEN_17954); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17956 = 8'h23 == cnt[7:0] ? $signed(32'she8bf) : $signed(_GEN_17955); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17957 = 8'h24 == cnt[7:0] ? $signed(32'she76c) : $signed(_GEN_17956); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17958 = 8'h25 == cnt[7:0] ? $signed(32'she610) : $signed(_GEN_17957); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17959 = 8'h26 == cnt[7:0] ? $signed(32'she4aa) : $signed(_GEN_17958); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17960 = 8'h27 == cnt[7:0] ? $signed(32'she33c) : $signed(_GEN_17959); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17961 = 8'h28 == cnt[7:0] ? $signed(32'she1c6) : $signed(_GEN_17960); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17962 = 8'h29 == cnt[7:0] ? $signed(32'she046) : $signed(_GEN_17961); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17963 = 8'h2a == cnt[7:0] ? $signed(32'shdebe) : $signed(_GEN_17962); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17964 = 8'h2b == cnt[7:0] ? $signed(32'shdd2d) : $signed(_GEN_17963); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17965 = 8'h2c == cnt[7:0] ? $signed(32'shdb94) : $signed(_GEN_17964); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17966 = 8'h2d == cnt[7:0] ? $signed(32'shd9f2) : $signed(_GEN_17965); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17967 = 8'h2e == cnt[7:0] ? $signed(32'shd848) : $signed(_GEN_17966); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17968 = 8'h2f == cnt[7:0] ? $signed(32'shd696) : $signed(_GEN_17967); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17969 = 8'h30 == cnt[7:0] ? $signed(32'shd4db) : $signed(_GEN_17968); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17970 = 8'h31 == cnt[7:0] ? $signed(32'shd318) : $signed(_GEN_17969); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17971 = 8'h32 == cnt[7:0] ? $signed(32'shd14d) : $signed(_GEN_17970); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17972 = 8'h33 == cnt[7:0] ? $signed(32'shcf7a) : $signed(_GEN_17971); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17973 = 8'h34 == cnt[7:0] ? $signed(32'shcd9f) : $signed(_GEN_17972); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17974 = 8'h35 == cnt[7:0] ? $signed(32'shcbbc) : $signed(_GEN_17973); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17975 = 8'h36 == cnt[7:0] ? $signed(32'shc9d1) : $signed(_GEN_17974); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17976 = 8'h37 == cnt[7:0] ? $signed(32'shc7de) : $signed(_GEN_17975); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17977 = 8'h38 == cnt[7:0] ? $signed(32'shc5e4) : $signed(_GEN_17976); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17978 = 8'h39 == cnt[7:0] ? $signed(32'shc3e2) : $signed(_GEN_17977); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17979 = 8'h3a == cnt[7:0] ? $signed(32'shc1d8) : $signed(_GEN_17978); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17980 = 8'h3b == cnt[7:0] ? $signed(32'shbfc7) : $signed(_GEN_17979); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17981 = 8'h3c == cnt[7:0] ? $signed(32'shbdaf) : $signed(_GEN_17980); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17982 = 8'h3d == cnt[7:0] ? $signed(32'shbb8f) : $signed(_GEN_17981); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17983 = 8'h3e == cnt[7:0] ? $signed(32'shb968) : $signed(_GEN_17982); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17984 = 8'h3f == cnt[7:0] ? $signed(32'shb73a) : $signed(_GEN_17983); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17985 = 8'h40 == cnt[7:0] ? $signed(32'shb505) : $signed(_GEN_17984); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17986 = 8'h41 == cnt[7:0] ? $signed(32'shb2c9) : $signed(_GEN_17985); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17987 = 8'h42 == cnt[7:0] ? $signed(32'shb086) : $signed(_GEN_17986); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17988 = 8'h43 == cnt[7:0] ? $signed(32'shae3c) : $signed(_GEN_17987); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17989 = 8'h44 == cnt[7:0] ? $signed(32'shabeb) : $signed(_GEN_17988); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17990 = 8'h45 == cnt[7:0] ? $signed(32'sha994) : $signed(_GEN_17989); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17991 = 8'h46 == cnt[7:0] ? $signed(32'sha736) : $signed(_GEN_17990); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17992 = 8'h47 == cnt[7:0] ? $signed(32'sha4d2) : $signed(_GEN_17991); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17993 = 8'h48 == cnt[7:0] ? $signed(32'sha268) : $signed(_GEN_17992); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17994 = 8'h49 == cnt[7:0] ? $signed(32'sh9ff7) : $signed(_GEN_17993); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17995 = 8'h4a == cnt[7:0] ? $signed(32'sh9d80) : $signed(_GEN_17994); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17996 = 8'h4b == cnt[7:0] ? $signed(32'sh9b03) : $signed(_GEN_17995); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17997 = 8'h4c == cnt[7:0] ? $signed(32'sh9880) : $signed(_GEN_17996); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17998 = 8'h4d == cnt[7:0] ? $signed(32'sh95f7) : $signed(_GEN_17997); // @[FFT.scala 34:12]
  wire [31:0] _GEN_17999 = 8'h4e == cnt[7:0] ? $signed(32'sh9368) : $signed(_GEN_17998); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18000 = 8'h4f == cnt[7:0] ? $signed(32'sh90d4) : $signed(_GEN_17999); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18001 = 8'h50 == cnt[7:0] ? $signed(32'sh8e3a) : $signed(_GEN_18000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18002 = 8'h51 == cnt[7:0] ? $signed(32'sh8b9a) : $signed(_GEN_18001); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18003 = 8'h52 == cnt[7:0] ? $signed(32'sh88f6) : $signed(_GEN_18002); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18004 = 8'h53 == cnt[7:0] ? $signed(32'sh864c) : $signed(_GEN_18003); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18005 = 8'h54 == cnt[7:0] ? $signed(32'sh839c) : $signed(_GEN_18004); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18006 = 8'h55 == cnt[7:0] ? $signed(32'sh80e8) : $signed(_GEN_18005); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18007 = 8'h56 == cnt[7:0] ? $signed(32'sh7e2f) : $signed(_GEN_18006); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18008 = 8'h57 == cnt[7:0] ? $signed(32'sh7b70) : $signed(_GEN_18007); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18009 = 8'h58 == cnt[7:0] ? $signed(32'sh78ad) : $signed(_GEN_18008); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18010 = 8'h59 == cnt[7:0] ? $signed(32'sh75e6) : $signed(_GEN_18009); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18011 = 8'h5a == cnt[7:0] ? $signed(32'sh731a) : $signed(_GEN_18010); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18012 = 8'h5b == cnt[7:0] ? $signed(32'sh7049) : $signed(_GEN_18011); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18013 = 8'h5c == cnt[7:0] ? $signed(32'sh6d74) : $signed(_GEN_18012); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18014 = 8'h5d == cnt[7:0] ? $signed(32'sh6a9b) : $signed(_GEN_18013); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18015 = 8'h5e == cnt[7:0] ? $signed(32'sh67be) : $signed(_GEN_18014); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18016 = 8'h5f == cnt[7:0] ? $signed(32'sh64dd) : $signed(_GEN_18015); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18017 = 8'h60 == cnt[7:0] ? $signed(32'sh61f8) : $signed(_GEN_18016); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18018 = 8'h61 == cnt[7:0] ? $signed(32'sh5f0f) : $signed(_GEN_18017); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18019 = 8'h62 == cnt[7:0] ? $signed(32'sh5c22) : $signed(_GEN_18018); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18020 = 8'h63 == cnt[7:0] ? $signed(32'sh5932) : $signed(_GEN_18019); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18021 = 8'h64 == cnt[7:0] ? $signed(32'sh563e) : $signed(_GEN_18020); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18022 = 8'h65 == cnt[7:0] ? $signed(32'sh5348) : $signed(_GEN_18021); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18023 = 8'h66 == cnt[7:0] ? $signed(32'sh504d) : $signed(_GEN_18022); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18024 = 8'h67 == cnt[7:0] ? $signed(32'sh4d50) : $signed(_GEN_18023); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18025 = 8'h68 == cnt[7:0] ? $signed(32'sh4a50) : $signed(_GEN_18024); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18026 = 8'h69 == cnt[7:0] ? $signed(32'sh474d) : $signed(_GEN_18025); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18027 = 8'h6a == cnt[7:0] ? $signed(32'sh4447) : $signed(_GEN_18026); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18028 = 8'h6b == cnt[7:0] ? $signed(32'sh413f) : $signed(_GEN_18027); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18029 = 8'h6c == cnt[7:0] ? $signed(32'sh3e34) : $signed(_GEN_18028); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18030 = 8'h6d == cnt[7:0] ? $signed(32'sh3b27) : $signed(_GEN_18029); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18031 = 8'h6e == cnt[7:0] ? $signed(32'sh3817) : $signed(_GEN_18030); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18032 = 8'h6f == cnt[7:0] ? $signed(32'sh3505) : $signed(_GEN_18031); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18033 = 8'h70 == cnt[7:0] ? $signed(32'sh31f1) : $signed(_GEN_18032); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18034 = 8'h71 == cnt[7:0] ? $signed(32'sh2edc) : $signed(_GEN_18033); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18035 = 8'h72 == cnt[7:0] ? $signed(32'sh2bc4) : $signed(_GEN_18034); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18036 = 8'h73 == cnt[7:0] ? $signed(32'sh28ab) : $signed(_GEN_18035); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18037 = 8'h74 == cnt[7:0] ? $signed(32'sh2590) : $signed(_GEN_18036); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18038 = 8'h75 == cnt[7:0] ? $signed(32'sh2274) : $signed(_GEN_18037); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18039 = 8'h76 == cnt[7:0] ? $signed(32'sh1f56) : $signed(_GEN_18038); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18040 = 8'h77 == cnt[7:0] ? $signed(32'sh1c38) : $signed(_GEN_18039); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18041 = 8'h78 == cnt[7:0] ? $signed(32'sh1918) : $signed(_GEN_18040); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18042 = 8'h79 == cnt[7:0] ? $signed(32'sh15f7) : $signed(_GEN_18041); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18043 = 8'h7a == cnt[7:0] ? $signed(32'sh12d5) : $signed(_GEN_18042); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18044 = 8'h7b == cnt[7:0] ? $signed(32'shfb3) : $signed(_GEN_18043); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18045 = 8'h7c == cnt[7:0] ? $signed(32'shc90) : $signed(_GEN_18044); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18046 = 8'h7d == cnt[7:0] ? $signed(32'sh96c) : $signed(_GEN_18045); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18047 = 8'h7e == cnt[7:0] ? $signed(32'sh648) : $signed(_GEN_18046); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18048 = 8'h7f == cnt[7:0] ? $signed(32'sh324) : $signed(_GEN_18047); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18049 = 8'h80 == cnt[7:0] ? $signed(32'sh0) : $signed(_GEN_18048); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18050 = 8'h81 == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_18049); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18051 = 8'h82 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_18050); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18052 = 8'h83 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_18051); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18053 = 8'h84 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_18052); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18054 = 8'h85 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_18053); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18055 = 8'h86 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_18054); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18056 = 8'h87 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_18055); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18057 = 8'h88 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_18056); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18058 = 8'h89 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_18057); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18059 = 8'h8a == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_18058); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18060 = 8'h8b == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_18059); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18061 = 8'h8c == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_18060); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18062 = 8'h8d == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_18061); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18063 = 8'h8e == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_18062); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18064 = 8'h8f == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_18063); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18065 = 8'h90 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_18064); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18066 = 8'h91 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_18065); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18067 = 8'h92 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_18066); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18068 = 8'h93 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_18067); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18069 = 8'h94 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_18068); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18070 = 8'h95 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_18069); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18071 = 8'h96 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_18070); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18072 = 8'h97 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_18071); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18073 = 8'h98 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_18072); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18074 = 8'h99 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_18073); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18075 = 8'h9a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_18074); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18076 = 8'h9b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_18075); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18077 = 8'h9c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_18076); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18078 = 8'h9d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_18077); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18079 = 8'h9e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_18078); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18080 = 8'h9f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_18079); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18081 = 8'ha0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_18080); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18082 = 8'ha1 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_18081); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18083 = 8'ha2 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_18082); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18084 = 8'ha3 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_18083); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18085 = 8'ha4 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_18084); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18086 = 8'ha5 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_18085); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18087 = 8'ha6 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_18086); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18088 = 8'ha7 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_18087); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18089 = 8'ha8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_18088); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18090 = 8'ha9 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_18089); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18091 = 8'haa == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_18090); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18092 = 8'hab == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_18091); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18093 = 8'hac == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_18092); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18094 = 8'had == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_18093); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18095 = 8'hae == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_18094); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18096 = 8'haf == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_18095); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18097 = 8'hb0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_18096); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18098 = 8'hb1 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_18097); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18099 = 8'hb2 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_18098); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18100 = 8'hb3 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_18099); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18101 = 8'hb4 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_18100); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18102 = 8'hb5 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_18101); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18103 = 8'hb6 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_18102); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18104 = 8'hb7 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_18103); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18105 = 8'hb8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_18104); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18106 = 8'hb9 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_18105); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18107 = 8'hba == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_18106); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18108 = 8'hbb == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_18107); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18109 = 8'hbc == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_18108); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18110 = 8'hbd == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_18109); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18111 = 8'hbe == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_18110); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18112 = 8'hbf == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_18111); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18113 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_18112); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18114 = 8'hc1 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_18113); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18115 = 8'hc2 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_18114); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18116 = 8'hc3 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_18115); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18117 = 8'hc4 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_18116); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18118 = 8'hc5 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_18117); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18119 = 8'hc6 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_18118); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18120 = 8'hc7 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_18119); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18121 = 8'hc8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_18120); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18122 = 8'hc9 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_18121); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18123 = 8'hca == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_18122); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18124 = 8'hcb == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_18123); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18125 = 8'hcc == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_18124); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18126 = 8'hcd == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_18125); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18127 = 8'hce == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_18126); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18128 = 8'hcf == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_18127); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18129 = 8'hd0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_18128); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18130 = 8'hd1 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_18129); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18131 = 8'hd2 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_18130); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18132 = 8'hd3 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_18131); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18133 = 8'hd4 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_18132); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18134 = 8'hd5 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_18133); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18135 = 8'hd6 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_18134); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18136 = 8'hd7 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_18135); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18137 = 8'hd8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_18136); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18138 = 8'hd9 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_18137); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18139 = 8'hda == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_18138); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18140 = 8'hdb == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_18139); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18141 = 8'hdc == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_18140); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18142 = 8'hdd == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_18141); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18143 = 8'hde == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_18142); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18144 = 8'hdf == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_18143); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18145 = 8'he0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_18144); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18146 = 8'he1 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_18145); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18147 = 8'he2 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_18146); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18148 = 8'he3 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_18147); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18149 = 8'he4 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_18148); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18150 = 8'he5 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_18149); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18151 = 8'he6 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_18150); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18152 = 8'he7 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_18151); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18153 = 8'he8 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_18152); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18154 = 8'he9 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_18153); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18155 = 8'hea == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_18154); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18156 = 8'heb == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_18155); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18157 = 8'hec == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_18156); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18158 = 8'hed == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_18157); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18159 = 8'hee == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_18158); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18160 = 8'hef == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_18159); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18161 = 8'hf0 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_18160); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18162 = 8'hf1 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_18161); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18163 = 8'hf2 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_18162); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18164 = 8'hf3 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_18163); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18165 = 8'hf4 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_18164); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18166 = 8'hf5 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_18165); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18167 = 8'hf6 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_18166); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18168 = 8'hf7 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_18167); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18169 = 8'hf8 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_18168); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18170 = 8'hf9 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_18169); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18171 = 8'hfa == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_18170); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18172 = 8'hfb == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_18171); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18173 = 8'hfc == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_18172); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18174 = 8'hfd == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_18173); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18175 = 8'hfe == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_18174); // @[FFT.scala 34:12]
  wire [31:0] _GEN_18178 = 8'h1 == cnt[7:0] ? $signed(-32'sh324) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18179 = 8'h2 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_18178); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18180 = 8'h3 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_18179); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18181 = 8'h4 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_18180); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18182 = 8'h5 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_18181); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18183 = 8'h6 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_18182); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18184 = 8'h7 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_18183); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18185 = 8'h8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_18184); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18186 = 8'h9 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_18185); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18187 = 8'ha == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_18186); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18188 = 8'hb == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_18187); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18189 = 8'hc == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_18188); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18190 = 8'hd == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_18189); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18191 = 8'he == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_18190); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18192 = 8'hf == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_18191); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18193 = 8'h10 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_18192); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18194 = 8'h11 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_18193); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18195 = 8'h12 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_18194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18196 = 8'h13 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_18195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18197 = 8'h14 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_18196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18198 = 8'h15 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_18197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18199 = 8'h16 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_18198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18200 = 8'h17 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_18199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18201 = 8'h18 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_18200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18202 = 8'h19 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_18201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18203 = 8'h1a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_18202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18204 = 8'h1b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_18203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18205 = 8'h1c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_18204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18206 = 8'h1d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_18205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18207 = 8'h1e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_18206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18208 = 8'h1f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_18207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18209 = 8'h20 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_18208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18210 = 8'h21 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_18209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18211 = 8'h22 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_18210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18212 = 8'h23 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_18211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18213 = 8'h24 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_18212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18214 = 8'h25 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_18213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18215 = 8'h26 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_18214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18216 = 8'h27 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_18215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18217 = 8'h28 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_18216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18218 = 8'h29 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_18217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18219 = 8'h2a == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_18218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18220 = 8'h2b == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_18219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18221 = 8'h2c == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_18220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18222 = 8'h2d == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_18221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18223 = 8'h2e == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_18222); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18224 = 8'h2f == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_18223); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18225 = 8'h30 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_18224); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18226 = 8'h31 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_18225); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18227 = 8'h32 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_18226); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18228 = 8'h33 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_18227); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18229 = 8'h34 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_18228); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18230 = 8'h35 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_18229); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18231 = 8'h36 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_18230); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18232 = 8'h37 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_18231); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18233 = 8'h38 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_18232); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18234 = 8'h39 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_18233); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18235 = 8'h3a == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_18234); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18236 = 8'h3b == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_18235); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18237 = 8'h3c == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_18236); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18238 = 8'h3d == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_18237); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18239 = 8'h3e == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_18238); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18240 = 8'h3f == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_18239); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18241 = 8'h40 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_18240); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18242 = 8'h41 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_18241); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18243 = 8'h42 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_18242); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18244 = 8'h43 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_18243); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18245 = 8'h44 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_18244); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18246 = 8'h45 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_18245); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18247 = 8'h46 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_18246); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18248 = 8'h47 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_18247); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18249 = 8'h48 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_18248); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18250 = 8'h49 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_18249); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18251 = 8'h4a == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_18250); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18252 = 8'h4b == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_18251); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18253 = 8'h4c == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_18252); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18254 = 8'h4d == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_18253); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18255 = 8'h4e == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_18254); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18256 = 8'h4f == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_18255); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18257 = 8'h50 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_18256); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18258 = 8'h51 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_18257); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18259 = 8'h52 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_18258); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18260 = 8'h53 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_18259); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18261 = 8'h54 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_18260); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18262 = 8'h55 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_18261); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18263 = 8'h56 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_18262); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18264 = 8'h57 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_18263); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18265 = 8'h58 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_18264); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18266 = 8'h59 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_18265); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18267 = 8'h5a == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_18266); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18268 = 8'h5b == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_18267); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18269 = 8'h5c == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_18268); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18270 = 8'h5d == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_18269); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18271 = 8'h5e == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_18270); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18272 = 8'h5f == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_18271); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18273 = 8'h60 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_18272); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18274 = 8'h61 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_18273); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18275 = 8'h62 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_18274); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18276 = 8'h63 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_18275); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18277 = 8'h64 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_18276); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18278 = 8'h65 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_18277); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18279 = 8'h66 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_18278); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18280 = 8'h67 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_18279); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18281 = 8'h68 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_18280); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18282 = 8'h69 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_18281); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18283 = 8'h6a == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_18282); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18284 = 8'h6b == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_18283); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18285 = 8'h6c == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_18284); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18286 = 8'h6d == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_18285); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18287 = 8'h6e == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_18286); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18288 = 8'h6f == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_18287); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18289 = 8'h70 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_18288); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18290 = 8'h71 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_18289); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18291 = 8'h72 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_18290); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18292 = 8'h73 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_18291); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18293 = 8'h74 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_18292); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18294 = 8'h75 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_18293); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18295 = 8'h76 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_18294); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18296 = 8'h77 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_18295); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18297 = 8'h78 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_18296); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18298 = 8'h79 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_18297); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18299 = 8'h7a == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_18298); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18300 = 8'h7b == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_18299); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18301 = 8'h7c == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_18300); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18302 = 8'h7d == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_18301); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18303 = 8'h7e == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_18302); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18304 = 8'h7f == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_18303); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18305 = 8'h80 == cnt[7:0] ? $signed(-32'sh10000) : $signed(_GEN_18304); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18306 = 8'h81 == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_18305); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18307 = 8'h82 == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_18306); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18308 = 8'h83 == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_18307); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18309 = 8'h84 == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_18308); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18310 = 8'h85 == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_18309); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18311 = 8'h86 == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_18310); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18312 = 8'h87 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_18311); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18313 = 8'h88 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_18312); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18314 = 8'h89 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_18313); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18315 = 8'h8a == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_18314); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18316 = 8'h8b == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_18315); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18317 = 8'h8c == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_18316); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18318 = 8'h8d == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_18317); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18319 = 8'h8e == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_18318); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18320 = 8'h8f == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_18319); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18321 = 8'h90 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_18320); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18322 = 8'h91 == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_18321); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18323 = 8'h92 == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_18322); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18324 = 8'h93 == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_18323); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18325 = 8'h94 == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_18324); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18326 = 8'h95 == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_18325); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18327 = 8'h96 == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_18326); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18328 = 8'h97 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_18327); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18329 = 8'h98 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_18328); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18330 = 8'h99 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_18329); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18331 = 8'h9a == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_18330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18332 = 8'h9b == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_18331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18333 = 8'h9c == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_18332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18334 = 8'h9d == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_18333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18335 = 8'h9e == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_18334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18336 = 8'h9f == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_18335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18337 = 8'ha0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_18336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18338 = 8'ha1 == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_18337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18339 = 8'ha2 == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_18338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18340 = 8'ha3 == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_18339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18341 = 8'ha4 == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_18340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18342 = 8'ha5 == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_18341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18343 = 8'ha6 == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_18342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18344 = 8'ha7 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_18343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18345 = 8'ha8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_18344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18346 = 8'ha9 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_18345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18347 = 8'haa == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_18346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18348 = 8'hab == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_18347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18349 = 8'hac == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_18348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18350 = 8'had == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_18349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18351 = 8'hae == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_18350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18352 = 8'haf == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_18351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18353 = 8'hb0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_18352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18354 = 8'hb1 == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_18353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18355 = 8'hb2 == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_18354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18356 = 8'hb3 == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_18355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18357 = 8'hb4 == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_18356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18358 = 8'hb5 == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_18357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18359 = 8'hb6 == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_18358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18360 = 8'hb7 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_18359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18361 = 8'hb8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_18360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18362 = 8'hb9 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_18361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18363 = 8'hba == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_18362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18364 = 8'hbb == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_18363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18365 = 8'hbc == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_18364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18366 = 8'hbd == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_18365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18367 = 8'hbe == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_18366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18368 = 8'hbf == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_18367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18369 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_18368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18370 = 8'hc1 == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_18369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18371 = 8'hc2 == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_18370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18372 = 8'hc3 == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_18371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18373 = 8'hc4 == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_18372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18374 = 8'hc5 == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_18373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18375 = 8'hc6 == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_18374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18376 = 8'hc7 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_18375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18377 = 8'hc8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_18376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18378 = 8'hc9 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_18377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18379 = 8'hca == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_18378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18380 = 8'hcb == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_18379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18381 = 8'hcc == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_18380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18382 = 8'hcd == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_18381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18383 = 8'hce == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_18382); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18384 = 8'hcf == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_18383); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18385 = 8'hd0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_18384); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18386 = 8'hd1 == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_18385); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18387 = 8'hd2 == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_18386); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18388 = 8'hd3 == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_18387); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18389 = 8'hd4 == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_18388); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18390 = 8'hd5 == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_18389); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18391 = 8'hd6 == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_18390); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18392 = 8'hd7 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_18391); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18393 = 8'hd8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_18392); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18394 = 8'hd9 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_18393); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18395 = 8'hda == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_18394); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18396 = 8'hdb == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_18395); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18397 = 8'hdc == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_18396); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18398 = 8'hdd == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_18397); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18399 = 8'hde == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_18398); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18400 = 8'hdf == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_18399); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18401 = 8'he0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_18400); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18402 = 8'he1 == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_18401); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18403 = 8'he2 == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_18402); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18404 = 8'he3 == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_18403); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18405 = 8'he4 == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_18404); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18406 = 8'he5 == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_18405); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18407 = 8'he6 == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_18406); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18408 = 8'he7 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_18407); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18409 = 8'he8 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_18408); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18410 = 8'he9 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_18409); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18411 = 8'hea == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_18410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18412 = 8'heb == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_18411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18413 = 8'hec == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_18412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18414 = 8'hed == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_18413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18415 = 8'hee == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_18414); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18416 = 8'hef == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_18415); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18417 = 8'hf0 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_18416); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18418 = 8'hf1 == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_18417); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18419 = 8'hf2 == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_18418); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18420 = 8'hf3 == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_18419); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18421 = 8'hf4 == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_18420); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18422 = 8'hf5 == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_18421); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18423 = 8'hf6 == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_18422); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18424 = 8'hf7 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_18423); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18425 = 8'hf8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_18424); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18426 = 8'hf9 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_18425); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18427 = 8'hfa == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_18426); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18428 = 8'hfb == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_18427); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18429 = 8'hfc == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_18428); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18430 = 8'hfd == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_18429); // @[FFT.scala 35:12]
  wire [31:0] _GEN_18431 = 8'hfe == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_18430); // @[FFT.scala 35:12]
  reg [31:0] _T_5586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10754;
  reg [31:0] _T_5586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10755;
  reg [31:0] _T_5587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10756;
  reg [31:0] _T_5587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10757;
  reg [31:0] _T_5588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10758;
  reg [31:0] _T_5588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10759;
  reg [31:0] _T_5589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10760;
  reg [31:0] _T_5589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10761;
  reg [31:0] _T_5590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10762;
  reg [31:0] _T_5590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10763;
  reg [31:0] _T_5591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10764;
  reg [31:0] _T_5591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10765;
  reg [31:0] _T_5592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10766;
  reg [31:0] _T_5592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10767;
  reg [31:0] _T_5593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10768;
  reg [31:0] _T_5593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10769;
  reg [31:0] _T_5594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10770;
  reg [31:0] _T_5594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10771;
  reg [31:0] _T_5595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10772;
  reg [31:0] _T_5595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10773;
  reg [31:0] _T_5596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10774;
  reg [31:0] _T_5596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10775;
  reg [31:0] _T_5597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10776;
  reg [31:0] _T_5597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10777;
  reg [31:0] _T_5598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10778;
  reg [31:0] _T_5598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10779;
  reg [31:0] _T_5599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10780;
  reg [31:0] _T_5599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10781;
  reg [31:0] _T_5600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10782;
  reg [31:0] _T_5600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10783;
  reg [31:0] _T_5601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10784;
  reg [31:0] _T_5601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10785;
  reg [31:0] _T_5602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10786;
  reg [31:0] _T_5602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10787;
  reg [31:0] _T_5603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10788;
  reg [31:0] _T_5603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10789;
  reg [31:0] _T_5604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10790;
  reg [31:0] _T_5604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10791;
  reg [31:0] _T_5605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10792;
  reg [31:0] _T_5605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10793;
  reg [31:0] _T_5606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10794;
  reg [31:0] _T_5606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10795;
  reg [31:0] _T_5607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10796;
  reg [31:0] _T_5607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10797;
  reg [31:0] _T_5608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10798;
  reg [31:0] _T_5608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10799;
  reg [31:0] _T_5609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10800;
  reg [31:0] _T_5609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10801;
  reg [31:0] _T_5610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10802;
  reg [31:0] _T_5610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10803;
  reg [31:0] _T_5611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10804;
  reg [31:0] _T_5611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10805;
  reg [31:0] _T_5612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10806;
  reg [31:0] _T_5612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10807;
  reg [31:0] _T_5613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10808;
  reg [31:0] _T_5613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10809;
  reg [31:0] _T_5614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10810;
  reg [31:0] _T_5614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10811;
  reg [31:0] _T_5615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10812;
  reg [31:0] _T_5615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10813;
  reg [31:0] _T_5616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10814;
  reg [31:0] _T_5616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10815;
  reg [31:0] _T_5617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10816;
  reg [31:0] _T_5617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10817;
  reg [31:0] _T_5618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10818;
  reg [31:0] _T_5618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10819;
  reg [31:0] _T_5619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10820;
  reg [31:0] _T_5619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10821;
  reg [31:0] _T_5620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10822;
  reg [31:0] _T_5620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10823;
  reg [31:0] _T_5621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10824;
  reg [31:0] _T_5621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10825;
  reg [31:0] _T_5622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10826;
  reg [31:0] _T_5622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10827;
  reg [31:0] _T_5623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10828;
  reg [31:0] _T_5623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10829;
  reg [31:0] _T_5624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10830;
  reg [31:0] _T_5624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10831;
  reg [31:0] _T_5625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10832;
  reg [31:0] _T_5625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10833;
  reg [31:0] _T_5626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10834;
  reg [31:0] _T_5626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10835;
  reg [31:0] _T_5627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10836;
  reg [31:0] _T_5627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10837;
  reg [31:0] _T_5628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10838;
  reg [31:0] _T_5628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10839;
  reg [31:0] _T_5629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10840;
  reg [31:0] _T_5629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10841;
  reg [31:0] _T_5630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10842;
  reg [31:0] _T_5630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10843;
  reg [31:0] _T_5631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10844;
  reg [31:0] _T_5631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10845;
  reg [31:0] _T_5632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10846;
  reg [31:0] _T_5632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10847;
  reg [31:0] _T_5633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10848;
  reg [31:0] _T_5633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10849;
  reg [31:0] _T_5634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10850;
  reg [31:0] _T_5634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10851;
  reg [31:0] _T_5635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10852;
  reg [31:0] _T_5635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10853;
  reg [31:0] _T_5636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10854;
  reg [31:0] _T_5636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10855;
  reg [31:0] _T_5637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10856;
  reg [31:0] _T_5637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10857;
  reg [31:0] _T_5638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10858;
  reg [31:0] _T_5638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10859;
  reg [31:0] _T_5639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10860;
  reg [31:0] _T_5639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10861;
  reg [31:0] _T_5640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10862;
  reg [31:0] _T_5640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10863;
  reg [31:0] _T_5641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10864;
  reg [31:0] _T_5641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10865;
  reg [31:0] _T_5642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10866;
  reg [31:0] _T_5642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10867;
  reg [31:0] _T_5643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10868;
  reg [31:0] _T_5643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10869;
  reg [31:0] _T_5644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10870;
  reg [31:0] _T_5644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10871;
  reg [31:0] _T_5645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10872;
  reg [31:0] _T_5645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10873;
  reg [31:0] _T_5646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10874;
  reg [31:0] _T_5646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10875;
  reg [31:0] _T_5647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10876;
  reg [31:0] _T_5647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10877;
  reg [31:0] _T_5648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10878;
  reg [31:0] _T_5648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10879;
  reg [31:0] _T_5649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10880;
  reg [31:0] _T_5649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10881;
  reg [31:0] _T_5650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10882;
  reg [31:0] _T_5650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10883;
  reg [31:0] _T_5651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10884;
  reg [31:0] _T_5651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10885;
  reg [31:0] _T_5652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10886;
  reg [31:0] _T_5652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10887;
  reg [31:0] _T_5653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10888;
  reg [31:0] _T_5653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10889;
  reg [31:0] _T_5654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10890;
  reg [31:0] _T_5654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10891;
  reg [31:0] _T_5655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10892;
  reg [31:0] _T_5655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10893;
  reg [31:0] _T_5656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10894;
  reg [31:0] _T_5656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10895;
  reg [31:0] _T_5657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10896;
  reg [31:0] _T_5657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10897;
  reg [31:0] _T_5658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10898;
  reg [31:0] _T_5658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10899;
  reg [31:0] _T_5659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10900;
  reg [31:0] _T_5659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10901;
  reg [31:0] _T_5660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10902;
  reg [31:0] _T_5660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10903;
  reg [31:0] _T_5661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10904;
  reg [31:0] _T_5661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10905;
  reg [31:0] _T_5662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10906;
  reg [31:0] _T_5662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10907;
  reg [31:0] _T_5663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10908;
  reg [31:0] _T_5663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10909;
  reg [31:0] _T_5664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10910;
  reg [31:0] _T_5664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10911;
  reg [31:0] _T_5665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10912;
  reg [31:0] _T_5665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10913;
  reg [31:0] _T_5666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10914;
  reg [31:0] _T_5666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10915;
  reg [31:0] _T_5667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10916;
  reg [31:0] _T_5667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10917;
  reg [31:0] _T_5668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10918;
  reg [31:0] _T_5668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10919;
  reg [31:0] _T_5669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10920;
  reg [31:0] _T_5669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10921;
  reg [31:0] _T_5670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10922;
  reg [31:0] _T_5670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10923;
  reg [31:0] _T_5671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10924;
  reg [31:0] _T_5671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10925;
  reg [31:0] _T_5672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10926;
  reg [31:0] _T_5672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10927;
  reg [31:0] _T_5673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10928;
  reg [31:0] _T_5673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10929;
  reg [31:0] _T_5674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10930;
  reg [31:0] _T_5674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10931;
  reg [31:0] _T_5675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10932;
  reg [31:0] _T_5675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10933;
  reg [31:0] _T_5676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10934;
  reg [31:0] _T_5676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10935;
  reg [31:0] _T_5677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10936;
  reg [31:0] _T_5677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10937;
  reg [31:0] _T_5678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10938;
  reg [31:0] _T_5678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10939;
  reg [31:0] _T_5679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10940;
  reg [31:0] _T_5679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10941;
  reg [31:0] _T_5680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10942;
  reg [31:0] _T_5680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10943;
  reg [31:0] _T_5681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10944;
  reg [31:0] _T_5681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10945;
  reg [31:0] _T_5682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10946;
  reg [31:0] _T_5682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10947;
  reg [31:0] _T_5683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10948;
  reg [31:0] _T_5683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10949;
  reg [31:0] _T_5684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10950;
  reg [31:0] _T_5684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10951;
  reg [31:0] _T_5685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10952;
  reg [31:0] _T_5685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10953;
  reg [31:0] _T_5686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10954;
  reg [31:0] _T_5686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10955;
  reg [31:0] _T_5687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10956;
  reg [31:0] _T_5687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10957;
  reg [31:0] _T_5688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10958;
  reg [31:0] _T_5688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10959;
  reg [31:0] _T_5689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10960;
  reg [31:0] _T_5689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10961;
  reg [31:0] _T_5690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10962;
  reg [31:0] _T_5690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10963;
  reg [31:0] _T_5691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10964;
  reg [31:0] _T_5691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10965;
  reg [31:0] _T_5692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10966;
  reg [31:0] _T_5692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10967;
  reg [31:0] _T_5693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10968;
  reg [31:0] _T_5693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10969;
  reg [31:0] _T_5694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10970;
  reg [31:0] _T_5694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10971;
  reg [31:0] _T_5695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10972;
  reg [31:0] _T_5695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10973;
  reg [31:0] _T_5696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10974;
  reg [31:0] _T_5696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10975;
  reg [31:0] _T_5697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10976;
  reg [31:0] _T_5697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10977;
  reg [31:0] _T_5698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10978;
  reg [31:0] _T_5698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10979;
  reg [31:0] _T_5699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10980;
  reg [31:0] _T_5699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10981;
  reg [31:0] _T_5700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10982;
  reg [31:0] _T_5700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10983;
  reg [31:0] _T_5701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10984;
  reg [31:0] _T_5701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10985;
  reg [31:0] _T_5702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10986;
  reg [31:0] _T_5702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10987;
  reg [31:0] _T_5703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10988;
  reg [31:0] _T_5703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10989;
  reg [31:0] _T_5704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10990;
  reg [31:0] _T_5704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10991;
  reg [31:0] _T_5705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10992;
  reg [31:0] _T_5705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10993;
  reg [31:0] _T_5706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10994;
  reg [31:0] _T_5706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10995;
  reg [31:0] _T_5707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10996;
  reg [31:0] _T_5707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10997;
  reg [31:0] _T_5708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10998;
  reg [31:0] _T_5708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10999;
  reg [31:0] _T_5709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11000;
  reg [31:0] _T_5709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11001;
  reg [31:0] _T_5710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11002;
  reg [31:0] _T_5710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11003;
  reg [31:0] _T_5711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11004;
  reg [31:0] _T_5711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11005;
  reg [31:0] _T_5712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11006;
  reg [31:0] _T_5712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11007;
  reg [31:0] _T_5713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11008;
  reg [31:0] _T_5713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11009;
  reg [31:0] _T_5714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11010;
  reg [31:0] _T_5714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11011;
  reg [31:0] _T_5715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11012;
  reg [31:0] _T_5715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11013;
  reg [31:0] _T_5716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11014;
  reg [31:0] _T_5716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11015;
  reg [31:0] _T_5717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11016;
  reg [31:0] _T_5717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11017;
  reg [31:0] _T_5718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11018;
  reg [31:0] _T_5718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11019;
  reg [31:0] _T_5719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11020;
  reg [31:0] _T_5719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11021;
  reg [31:0] _T_5720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11022;
  reg [31:0] _T_5720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11023;
  reg [31:0] _T_5721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11024;
  reg [31:0] _T_5721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11025;
  reg [31:0] _T_5722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11026;
  reg [31:0] _T_5722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11027;
  reg [31:0] _T_5723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11028;
  reg [31:0] _T_5723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11029;
  reg [31:0] _T_5724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11030;
  reg [31:0] _T_5724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11031;
  reg [31:0] _T_5725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11032;
  reg [31:0] _T_5725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11033;
  reg [31:0] _T_5726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11034;
  reg [31:0] _T_5726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11035;
  reg [31:0] _T_5727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11036;
  reg [31:0] _T_5727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11037;
  reg [31:0] _T_5728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11038;
  reg [31:0] _T_5728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11039;
  reg [31:0] _T_5729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11040;
  reg [31:0] _T_5729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11041;
  reg [31:0] _T_5730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11042;
  reg [31:0] _T_5730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11043;
  reg [31:0] _T_5731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11044;
  reg [31:0] _T_5731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11045;
  reg [31:0] _T_5732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11046;
  reg [31:0] _T_5732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11047;
  reg [31:0] _T_5733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11048;
  reg [31:0] _T_5733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11049;
  reg [31:0] _T_5734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11050;
  reg [31:0] _T_5734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11051;
  reg [31:0] _T_5735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11052;
  reg [31:0] _T_5735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11053;
  reg [31:0] _T_5736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11054;
  reg [31:0] _T_5736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11055;
  reg [31:0] _T_5737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11056;
  reg [31:0] _T_5737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11057;
  reg [31:0] _T_5738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11058;
  reg [31:0] _T_5738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11059;
  reg [31:0] _T_5739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11060;
  reg [31:0] _T_5739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11061;
  reg [31:0] _T_5740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11062;
  reg [31:0] _T_5740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11063;
  reg [31:0] _T_5741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11064;
  reg [31:0] _T_5741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11065;
  reg [31:0] _T_5742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11066;
  reg [31:0] _T_5742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11067;
  reg [31:0] _T_5743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11068;
  reg [31:0] _T_5743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11069;
  reg [31:0] _T_5744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11070;
  reg [31:0] _T_5744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11071;
  reg [31:0] _T_5745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11072;
  reg [31:0] _T_5745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11073;
  reg [31:0] _T_5746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11074;
  reg [31:0] _T_5746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11075;
  reg [31:0] _T_5747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11076;
  reg [31:0] _T_5747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11077;
  reg [31:0] _T_5748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11078;
  reg [31:0] _T_5748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11079;
  reg [31:0] _T_5749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11080;
  reg [31:0] _T_5749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11081;
  reg [31:0] _T_5750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11082;
  reg [31:0] _T_5750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11083;
  reg [31:0] _T_5751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11084;
  reg [31:0] _T_5751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11085;
  reg [31:0] _T_5752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11086;
  reg [31:0] _T_5752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11087;
  reg [31:0] _T_5753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11088;
  reg [31:0] _T_5753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11089;
  reg [31:0] _T_5754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11090;
  reg [31:0] _T_5754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11091;
  reg [31:0] _T_5755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11092;
  reg [31:0] _T_5755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11093;
  reg [31:0] _T_5756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11094;
  reg [31:0] _T_5756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11095;
  reg [31:0] _T_5757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11096;
  reg [31:0] _T_5757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11097;
  reg [31:0] _T_5758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11098;
  reg [31:0] _T_5758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11099;
  reg [31:0] _T_5759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11100;
  reg [31:0] _T_5759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11101;
  reg [31:0] _T_5760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11102;
  reg [31:0] _T_5760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11103;
  reg [31:0] _T_5761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11104;
  reg [31:0] _T_5761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11105;
  reg [31:0] _T_5762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11106;
  reg [31:0] _T_5762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11107;
  reg [31:0] _T_5763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11108;
  reg [31:0] _T_5763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11109;
  reg [31:0] _T_5764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11110;
  reg [31:0] _T_5764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11111;
  reg [31:0] _T_5765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11112;
  reg [31:0] _T_5765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11113;
  reg [31:0] _T_5766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11114;
  reg [31:0] _T_5766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11115;
  reg [31:0] _T_5767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11116;
  reg [31:0] _T_5767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11117;
  reg [31:0] _T_5768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11118;
  reg [31:0] _T_5768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11119;
  reg [31:0] _T_5769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11120;
  reg [31:0] _T_5769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11121;
  reg [31:0] _T_5770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11122;
  reg [31:0] _T_5770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11123;
  reg [31:0] _T_5771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11124;
  reg [31:0] _T_5771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11125;
  reg [31:0] _T_5772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11126;
  reg [31:0] _T_5772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11127;
  reg [31:0] _T_5773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11128;
  reg [31:0] _T_5773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11129;
  reg [31:0] _T_5774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11130;
  reg [31:0] _T_5774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11131;
  reg [31:0] _T_5775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11132;
  reg [31:0] _T_5775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11133;
  reg [31:0] _T_5776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11134;
  reg [31:0] _T_5776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11135;
  reg [31:0] _T_5777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11136;
  reg [31:0] _T_5777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11137;
  reg [31:0] _T_5778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11138;
  reg [31:0] _T_5778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11139;
  reg [31:0] _T_5779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11140;
  reg [31:0] _T_5779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11141;
  reg [31:0] _T_5780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11142;
  reg [31:0] _T_5780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11143;
  reg [31:0] _T_5781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11144;
  reg [31:0] _T_5781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11145;
  reg [31:0] _T_5782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11146;
  reg [31:0] _T_5782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11147;
  reg [31:0] _T_5783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11148;
  reg [31:0] _T_5783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11149;
  reg [31:0] _T_5784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11150;
  reg [31:0] _T_5784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11151;
  reg [31:0] _T_5785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11152;
  reg [31:0] _T_5785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11153;
  reg [31:0] _T_5786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11154;
  reg [31:0] _T_5786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11155;
  reg [31:0] _T_5787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11156;
  reg [31:0] _T_5787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11157;
  reg [31:0] _T_5788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11158;
  reg [31:0] _T_5788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11159;
  reg [31:0] _T_5789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11160;
  reg [31:0] _T_5789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11161;
  reg [31:0] _T_5790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11162;
  reg [31:0] _T_5790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11163;
  reg [31:0] _T_5791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11164;
  reg [31:0] _T_5791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11165;
  reg [31:0] _T_5792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11166;
  reg [31:0] _T_5792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11167;
  reg [31:0] _T_5793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11168;
  reg [31:0] _T_5793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11169;
  reg [31:0] _T_5794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11170;
  reg [31:0] _T_5794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11171;
  reg [31:0] _T_5795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11172;
  reg [31:0] _T_5795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11173;
  reg [31:0] _T_5796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11174;
  reg [31:0] _T_5796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11175;
  reg [31:0] _T_5797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11176;
  reg [31:0] _T_5797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11177;
  reg [31:0] _T_5798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11178;
  reg [31:0] _T_5798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11179;
  reg [31:0] _T_5799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11180;
  reg [31:0] _T_5799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11181;
  reg [31:0] _T_5800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11182;
  reg [31:0] _T_5800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11183;
  reg [31:0] _T_5801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11184;
  reg [31:0] _T_5801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11185;
  reg [31:0] _T_5802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11186;
  reg [31:0] _T_5802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11187;
  reg [31:0] _T_5803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11188;
  reg [31:0] _T_5803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11189;
  reg [31:0] _T_5804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11190;
  reg [31:0] _T_5804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11191;
  reg [31:0] _T_5805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11192;
  reg [31:0] _T_5805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11193;
  reg [31:0] _T_5806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11194;
  reg [31:0] _T_5806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11195;
  reg [31:0] _T_5807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11196;
  reg [31:0] _T_5807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11197;
  reg [31:0] _T_5808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11198;
  reg [31:0] _T_5808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11199;
  reg [31:0] _T_5809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11200;
  reg [31:0] _T_5809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11201;
  reg [31:0] _T_5810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11202;
  reg [31:0] _T_5810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11203;
  reg [31:0] _T_5811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11204;
  reg [31:0] _T_5811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11205;
  reg [31:0] _T_5812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11206;
  reg [31:0] _T_5812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11207;
  reg [31:0] _T_5813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11208;
  reg [31:0] _T_5813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11209;
  reg [31:0] _T_5814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11210;
  reg [31:0] _T_5814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11211;
  reg [31:0] _T_5815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11212;
  reg [31:0] _T_5815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11213;
  reg [31:0] _T_5816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11214;
  reg [31:0] _T_5816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11215;
  reg [31:0] _T_5817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11216;
  reg [31:0] _T_5817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11217;
  reg [31:0] _T_5818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11218;
  reg [31:0] _T_5818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11219;
  reg [31:0] _T_5819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11220;
  reg [31:0] _T_5819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11221;
  reg [31:0] _T_5820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11222;
  reg [31:0] _T_5820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11223;
  reg [31:0] _T_5821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11224;
  reg [31:0] _T_5821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11225;
  reg [31:0] _T_5822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11226;
  reg [31:0] _T_5822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11227;
  reg [31:0] _T_5823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11228;
  reg [31:0] _T_5823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11229;
  reg [31:0] _T_5824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11230;
  reg [31:0] _T_5824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11231;
  reg [31:0] _T_5825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11232;
  reg [31:0] _T_5825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11233;
  reg [31:0] _T_5826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11234;
  reg [31:0] _T_5826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11235;
  reg [31:0] _T_5827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11236;
  reg [31:0] _T_5827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11237;
  reg [31:0] _T_5828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11238;
  reg [31:0] _T_5828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11239;
  reg [31:0] _T_5829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11240;
  reg [31:0] _T_5829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11241;
  reg [31:0] _T_5830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11242;
  reg [31:0] _T_5830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11243;
  reg [31:0] _T_5831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11244;
  reg [31:0] _T_5831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11245;
  reg [31:0] _T_5832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11246;
  reg [31:0] _T_5832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11247;
  reg [31:0] _T_5833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11248;
  reg [31:0] _T_5833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11249;
  reg [31:0] _T_5834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11250;
  reg [31:0] _T_5834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11251;
  reg [31:0] _T_5835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11252;
  reg [31:0] _T_5835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11253;
  reg [31:0] _T_5836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11254;
  reg [31:0] _T_5836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11255;
  reg [31:0] _T_5837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11256;
  reg [31:0] _T_5837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11257;
  reg [31:0] _T_5838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11258;
  reg [31:0] _T_5838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11259;
  reg [31:0] _T_5839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11260;
  reg [31:0] _T_5839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11261;
  reg [31:0] _T_5840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11262;
  reg [31:0] _T_5840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11263;
  reg [31:0] _T_5841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11264;
  reg [31:0] _T_5841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11265;
  reg [31:0] _T_5844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11266;
  reg [31:0] _T_5844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11267;
  reg [31:0] _T_5845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11268;
  reg [31:0] _T_5845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11269;
  reg [31:0] _T_5846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11270;
  reg [31:0] _T_5846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11271;
  reg [31:0] _T_5847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11272;
  reg [31:0] _T_5847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11273;
  reg [31:0] _T_5848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11274;
  reg [31:0] _T_5848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11275;
  reg [31:0] _T_5849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11276;
  reg [31:0] _T_5849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11277;
  reg [31:0] _T_5850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11278;
  reg [31:0] _T_5850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11279;
  reg [31:0] _T_5851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11280;
  reg [31:0] _T_5851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11281;
  reg [31:0] _T_5852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11282;
  reg [31:0] _T_5852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11283;
  reg [31:0] _T_5853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11284;
  reg [31:0] _T_5853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11285;
  reg [31:0] _T_5854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11286;
  reg [31:0] _T_5854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11287;
  reg [31:0] _T_5855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11288;
  reg [31:0] _T_5855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11289;
  reg [31:0] _T_5856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11290;
  reg [31:0] _T_5856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11291;
  reg [31:0] _T_5857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11292;
  reg [31:0] _T_5857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11293;
  reg [31:0] _T_5858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11294;
  reg [31:0] _T_5858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11295;
  reg [31:0] _T_5859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11296;
  reg [31:0] _T_5859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11297;
  reg [31:0] _T_5860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11298;
  reg [31:0] _T_5860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11299;
  reg [31:0] _T_5861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11300;
  reg [31:0] _T_5861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11301;
  reg [31:0] _T_5862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11302;
  reg [31:0] _T_5862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11303;
  reg [31:0] _T_5863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11304;
  reg [31:0] _T_5863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11305;
  reg [31:0] _T_5864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11306;
  reg [31:0] _T_5864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11307;
  reg [31:0] _T_5865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11308;
  reg [31:0] _T_5865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11309;
  reg [31:0] _T_5866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11310;
  reg [31:0] _T_5866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11311;
  reg [31:0] _T_5867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11312;
  reg [31:0] _T_5867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11313;
  reg [31:0] _T_5868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11314;
  reg [31:0] _T_5868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11315;
  reg [31:0] _T_5869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11316;
  reg [31:0] _T_5869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11317;
  reg [31:0] _T_5870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11318;
  reg [31:0] _T_5870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11319;
  reg [31:0] _T_5871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11320;
  reg [31:0] _T_5871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11321;
  reg [31:0] _T_5872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11322;
  reg [31:0] _T_5872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11323;
  reg [31:0] _T_5873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11324;
  reg [31:0] _T_5873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11325;
  reg [31:0] _T_5874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11326;
  reg [31:0] _T_5874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11327;
  reg [31:0] _T_5875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11328;
  reg [31:0] _T_5875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11329;
  reg [31:0] _T_5876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11330;
  reg [31:0] _T_5876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11331;
  reg [31:0] _T_5877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11332;
  reg [31:0] _T_5877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11333;
  reg [31:0] _T_5878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11334;
  reg [31:0] _T_5878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11335;
  reg [31:0] _T_5879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11336;
  reg [31:0] _T_5879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11337;
  reg [31:0] _T_5880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11338;
  reg [31:0] _T_5880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11339;
  reg [31:0] _T_5881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11340;
  reg [31:0] _T_5881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11341;
  reg [31:0] _T_5882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11342;
  reg [31:0] _T_5882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11343;
  reg [31:0] _T_5883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11344;
  reg [31:0] _T_5883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11345;
  reg [31:0] _T_5884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11346;
  reg [31:0] _T_5884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11347;
  reg [31:0] _T_5885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11348;
  reg [31:0] _T_5885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11349;
  reg [31:0] _T_5886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11350;
  reg [31:0] _T_5886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11351;
  reg [31:0] _T_5887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11352;
  reg [31:0] _T_5887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11353;
  reg [31:0] _T_5888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11354;
  reg [31:0] _T_5888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11355;
  reg [31:0] _T_5889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11356;
  reg [31:0] _T_5889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11357;
  reg [31:0] _T_5890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11358;
  reg [31:0] _T_5890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11359;
  reg [31:0] _T_5891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11360;
  reg [31:0] _T_5891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11361;
  reg [31:0] _T_5892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11362;
  reg [31:0] _T_5892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11363;
  reg [31:0] _T_5893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11364;
  reg [31:0] _T_5893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11365;
  reg [31:0] _T_5894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11366;
  reg [31:0] _T_5894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11367;
  reg [31:0] _T_5895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11368;
  reg [31:0] _T_5895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11369;
  reg [31:0] _T_5896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11370;
  reg [31:0] _T_5896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11371;
  reg [31:0] _T_5897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11372;
  reg [31:0] _T_5897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11373;
  reg [31:0] _T_5898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11374;
  reg [31:0] _T_5898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11375;
  reg [31:0] _T_5899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11376;
  reg [31:0] _T_5899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11377;
  reg [31:0] _T_5900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11378;
  reg [31:0] _T_5900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11379;
  reg [31:0] _T_5901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11380;
  reg [31:0] _T_5901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11381;
  reg [31:0] _T_5902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11382;
  reg [31:0] _T_5902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11383;
  reg [31:0] _T_5903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11384;
  reg [31:0] _T_5903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11385;
  reg [31:0] _T_5904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11386;
  reg [31:0] _T_5904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11387;
  reg [31:0] _T_5905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11388;
  reg [31:0] _T_5905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11389;
  reg [31:0] _T_5906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11390;
  reg [31:0] _T_5906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11391;
  reg [31:0] _T_5907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11392;
  reg [31:0] _T_5907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11393;
  reg [31:0] _T_5908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11394;
  reg [31:0] _T_5908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11395;
  reg [31:0] _T_5909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11396;
  reg [31:0] _T_5909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11397;
  reg [31:0] _T_5910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11398;
  reg [31:0] _T_5910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11399;
  reg [31:0] _T_5911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11400;
  reg [31:0] _T_5911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11401;
  reg [31:0] _T_5912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11402;
  reg [31:0] _T_5912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11403;
  reg [31:0] _T_5913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11404;
  reg [31:0] _T_5913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11405;
  reg [31:0] _T_5914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11406;
  reg [31:0] _T_5914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11407;
  reg [31:0] _T_5915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11408;
  reg [31:0] _T_5915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11409;
  reg [31:0] _T_5916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11410;
  reg [31:0] _T_5916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11411;
  reg [31:0] _T_5917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11412;
  reg [31:0] _T_5917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11413;
  reg [31:0] _T_5918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11414;
  reg [31:0] _T_5918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11415;
  reg [31:0] _T_5919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11416;
  reg [31:0] _T_5919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11417;
  reg [31:0] _T_5920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11418;
  reg [31:0] _T_5920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11419;
  reg [31:0] _T_5921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11420;
  reg [31:0] _T_5921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11421;
  reg [31:0] _T_5922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11422;
  reg [31:0] _T_5922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11423;
  reg [31:0] _T_5923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11424;
  reg [31:0] _T_5923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11425;
  reg [31:0] _T_5924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11426;
  reg [31:0] _T_5924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11427;
  reg [31:0] _T_5925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11428;
  reg [31:0] _T_5925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11429;
  reg [31:0] _T_5926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11430;
  reg [31:0] _T_5926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11431;
  reg [31:0] _T_5927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11432;
  reg [31:0] _T_5927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11433;
  reg [31:0] _T_5928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11434;
  reg [31:0] _T_5928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11435;
  reg [31:0] _T_5929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11436;
  reg [31:0] _T_5929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11437;
  reg [31:0] _T_5930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11438;
  reg [31:0] _T_5930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11439;
  reg [31:0] _T_5931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11440;
  reg [31:0] _T_5931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11441;
  reg [31:0] _T_5932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11442;
  reg [31:0] _T_5932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11443;
  reg [31:0] _T_5933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11444;
  reg [31:0] _T_5933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11445;
  reg [31:0] _T_5934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11446;
  reg [31:0] _T_5934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11447;
  reg [31:0] _T_5935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11448;
  reg [31:0] _T_5935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11449;
  reg [31:0] _T_5936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11450;
  reg [31:0] _T_5936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11451;
  reg [31:0] _T_5937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11452;
  reg [31:0] _T_5937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11453;
  reg [31:0] _T_5938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11454;
  reg [31:0] _T_5938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11455;
  reg [31:0] _T_5939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11456;
  reg [31:0] _T_5939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11457;
  reg [31:0] _T_5940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11458;
  reg [31:0] _T_5940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11459;
  reg [31:0] _T_5941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11460;
  reg [31:0] _T_5941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11461;
  reg [31:0] _T_5942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11462;
  reg [31:0] _T_5942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11463;
  reg [31:0] _T_5943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11464;
  reg [31:0] _T_5943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11465;
  reg [31:0] _T_5944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11466;
  reg [31:0] _T_5944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11467;
  reg [31:0] _T_5945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11468;
  reg [31:0] _T_5945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11469;
  reg [31:0] _T_5946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11470;
  reg [31:0] _T_5946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11471;
  reg [31:0] _T_5947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11472;
  reg [31:0] _T_5947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11473;
  reg [31:0] _T_5948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11474;
  reg [31:0] _T_5948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11475;
  reg [31:0] _T_5949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11476;
  reg [31:0] _T_5949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11477;
  reg [31:0] _T_5950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11478;
  reg [31:0] _T_5950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11479;
  reg [31:0] _T_5951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11480;
  reg [31:0] _T_5951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11481;
  reg [31:0] _T_5952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11482;
  reg [31:0] _T_5952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11483;
  reg [31:0] _T_5953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11484;
  reg [31:0] _T_5953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11485;
  reg [31:0] _T_5954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11486;
  reg [31:0] _T_5954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11487;
  reg [31:0] _T_5955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11488;
  reg [31:0] _T_5955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11489;
  reg [31:0] _T_5956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11490;
  reg [31:0] _T_5956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11491;
  reg [31:0] _T_5957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11492;
  reg [31:0] _T_5957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11493;
  reg [31:0] _T_5958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11494;
  reg [31:0] _T_5958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11495;
  reg [31:0] _T_5959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11496;
  reg [31:0] _T_5959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11497;
  reg [31:0] _T_5960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11498;
  reg [31:0] _T_5960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11499;
  reg [31:0] _T_5961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11500;
  reg [31:0] _T_5961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11501;
  reg [31:0] _T_5962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11502;
  reg [31:0] _T_5962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11503;
  reg [31:0] _T_5963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11504;
  reg [31:0] _T_5963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11505;
  reg [31:0] _T_5964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11506;
  reg [31:0] _T_5964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11507;
  reg [31:0] _T_5965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11508;
  reg [31:0] _T_5965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11509;
  reg [31:0] _T_5966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11510;
  reg [31:0] _T_5966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11511;
  reg [31:0] _T_5967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11512;
  reg [31:0] _T_5967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11513;
  reg [31:0] _T_5968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11514;
  reg [31:0] _T_5968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11515;
  reg [31:0] _T_5969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11516;
  reg [31:0] _T_5969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11517;
  reg [31:0] _T_5970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11518;
  reg [31:0] _T_5970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11519;
  reg [31:0] _T_5971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11520;
  reg [31:0] _T_5971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11521;
  wire [31:0] _GEN_19202 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19203 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_19202); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19204 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_19203); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19205 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_19204); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19206 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_19205); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19207 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_19206); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19208 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_19207); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19209 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_19208); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19210 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_19209); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19211 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_19210); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19212 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_19211); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19213 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_19212); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19214 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_19213); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19215 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_19214); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19216 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_19215); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19217 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_19216); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19218 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_19217); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19219 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_19218); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19220 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_19219); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19221 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_19220); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19222 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_19221); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19223 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_19222); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19224 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_19223); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19225 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_19224); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19226 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_19225); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19227 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_19226); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19228 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_19227); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19229 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_19228); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19230 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_19229); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19231 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_19230); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19232 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_19231); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19233 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_19232); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19234 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_19233); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19235 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_19234); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19236 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_19235); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19237 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_19236); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19238 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_19237); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19239 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_19238); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19240 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_19239); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19241 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_19240); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19242 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_19241); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19243 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_19242); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19244 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_19243); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19245 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_19244); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19246 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_19245); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19247 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_19246); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19248 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_19247); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19249 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_19248); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19250 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_19249); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19251 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_19250); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19252 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_19251); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19253 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_19252); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19254 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_19253); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19255 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_19254); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19256 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_19255); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19257 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_19256); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19258 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_19257); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19259 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_19258); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19260 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_19259); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19261 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_19260); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19262 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_19261); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19263 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_19262); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19264 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_19263); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19265 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_19264); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19266 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_19265); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19267 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_19266); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19268 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_19267); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19269 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_19268); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19270 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_19269); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19271 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_19270); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19272 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_19271); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19273 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_19272); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19274 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_19273); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19275 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_19274); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19276 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_19275); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19277 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_19276); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19278 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_19277); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19279 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_19278); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19280 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_19279); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19281 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_19280); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19282 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_19281); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19283 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_19282); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19284 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_19283); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19285 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_19284); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19286 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_19285); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19287 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_19286); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19288 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_19287); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19289 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19288); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19290 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_19289); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19291 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_19290); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19292 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_19291); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19293 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_19292); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19294 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_19293); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19295 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_19294); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19296 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_19295); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19297 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_19296); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19298 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_19297); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19299 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_19298); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19300 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_19299); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19301 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_19300); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19302 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_19301); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19303 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_19302); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19304 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_19303); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19305 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_19304); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19306 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_19305); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19307 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_19306); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19308 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_19307); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19309 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_19308); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19310 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_19309); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19311 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_19310); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19312 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_19311); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19313 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_19312); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19314 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_19313); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19315 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_19314); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19316 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_19315); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19317 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_19316); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19318 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_19317); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19319 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_19318); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19320 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_19319); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19321 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_19320); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19322 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_19321); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19323 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_19322); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19324 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_19323); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19325 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_19324); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19326 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_19325); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19327 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_19326); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19330 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19331 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_19330); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19332 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_19331); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19333 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_19332); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19334 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_19333); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19335 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_19334); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19336 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_19335); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19337 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_19336); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19338 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_19337); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19339 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_19338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19340 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_19339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19341 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_19340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19342 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_19341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19343 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_19342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19344 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_19343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19345 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_19344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19346 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_19345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19347 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_19346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19348 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_19347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19349 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_19348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19350 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_19349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19351 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_19350); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19352 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_19351); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19353 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19352); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19354 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_19353); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19355 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_19354); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19356 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_19355); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19357 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_19356); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19358 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_19357); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19359 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_19358); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19360 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_19359); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19361 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_19360); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19362 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_19361); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19363 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_19362); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19364 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_19363); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19365 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_19364); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19366 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_19365); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19367 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_19366); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19368 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_19367); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19369 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_19368); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19370 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_19369); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19371 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_19370); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19372 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_19371); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19373 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_19372); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19374 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_19373); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19375 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_19374); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19376 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_19375); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19377 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_19376); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19378 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_19377); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19379 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_19378); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19380 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_19379); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19381 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_19380); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19382 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_19381); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19383 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_19382); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19384 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_19383); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19385 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_19384); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19386 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_19385); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19387 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_19386); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19388 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_19387); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19389 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_19388); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19390 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_19389); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19391 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_19390); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19392 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_19391); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19393 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_19392); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19394 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_19393); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19395 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_19394); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19396 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_19395); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19397 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_19396); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19398 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_19397); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19399 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_19398); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19400 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_19399); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19401 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_19400); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19402 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_19401); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19403 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_19402); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19404 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_19403); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19405 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_19404); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19406 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_19405); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19407 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_19406); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19408 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_19407); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19409 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_19408); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19410 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_19409); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19411 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_19410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19412 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_19411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19413 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_19412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19414 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_19413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19415 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_19414); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19416 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_19415); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19417 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_19416); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19418 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_19417); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19419 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_19418); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19420 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_19419); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19421 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_19420); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19422 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_19421); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19423 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_19422); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19424 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_19423); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19425 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_19424); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19426 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_19425); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19427 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_19426); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19428 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_19427); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19429 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_19428); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19430 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_19429); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19431 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_19430); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19432 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_19431); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19433 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19432); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19434 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_19433); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19435 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_19434); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19436 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_19435); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19437 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_19436); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19438 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_19437); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19439 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_19438); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19440 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_19439); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19441 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_19440); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19442 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_19441); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19443 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_19442); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19444 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_19443); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19445 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_19444); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19446 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_19445); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19447 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_19446); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19448 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_19447); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19449 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_19448); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19450 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_19449); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19451 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_19450); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19452 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_19451); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19453 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_19452); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19454 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_19453); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19455 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_19454); // @[FFT.scala 35:12]
  reg [31:0] _T_5977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11522;
  reg [31:0] _T_5977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11523;
  reg [31:0] _T_5978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11524;
  reg [31:0] _T_5978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11525;
  reg [31:0] _T_5979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11526;
  reg [31:0] _T_5979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11527;
  reg [31:0] _T_5980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11528;
  reg [31:0] _T_5980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11529;
  reg [31:0] _T_5981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11530;
  reg [31:0] _T_5981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11531;
  reg [31:0] _T_5982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11532;
  reg [31:0] _T_5982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11533;
  reg [31:0] _T_5983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11534;
  reg [31:0] _T_5983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11535;
  reg [31:0] _T_5984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11536;
  reg [31:0] _T_5984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11537;
  reg [31:0] _T_5985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11538;
  reg [31:0] _T_5985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11539;
  reg [31:0] _T_5986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11540;
  reg [31:0] _T_5986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11541;
  reg [31:0] _T_5987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11542;
  reg [31:0] _T_5987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11543;
  reg [31:0] _T_5988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11544;
  reg [31:0] _T_5988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11545;
  reg [31:0] _T_5989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11546;
  reg [31:0] _T_5989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11547;
  reg [31:0] _T_5990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11548;
  reg [31:0] _T_5990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11549;
  reg [31:0] _T_5991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11550;
  reg [31:0] _T_5991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11551;
  reg [31:0] _T_5992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11552;
  reg [31:0] _T_5992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11553;
  reg [31:0] _T_5993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11554;
  reg [31:0] _T_5993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11555;
  reg [31:0] _T_5994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11556;
  reg [31:0] _T_5994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11557;
  reg [31:0] _T_5995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11558;
  reg [31:0] _T_5995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11559;
  reg [31:0] _T_5996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11560;
  reg [31:0] _T_5996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11561;
  reg [31:0] _T_5997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11562;
  reg [31:0] _T_5997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11563;
  reg [31:0] _T_5998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11564;
  reg [31:0] _T_5998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11565;
  reg [31:0] _T_5999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11566;
  reg [31:0] _T_5999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11567;
  reg [31:0] _T_6000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11568;
  reg [31:0] _T_6000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11569;
  reg [31:0] _T_6001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11570;
  reg [31:0] _T_6001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11571;
  reg [31:0] _T_6002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11572;
  reg [31:0] _T_6002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11573;
  reg [31:0] _T_6003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11574;
  reg [31:0] _T_6003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11575;
  reg [31:0] _T_6004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11576;
  reg [31:0] _T_6004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11577;
  reg [31:0] _T_6005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11578;
  reg [31:0] _T_6005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11579;
  reg [31:0] _T_6006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11580;
  reg [31:0] _T_6006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11581;
  reg [31:0] _T_6007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11582;
  reg [31:0] _T_6007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11583;
  reg [31:0] _T_6008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11584;
  reg [31:0] _T_6008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11585;
  reg [31:0] _T_6009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11586;
  reg [31:0] _T_6009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11587;
  reg [31:0] _T_6010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11588;
  reg [31:0] _T_6010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11589;
  reg [31:0] _T_6011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11590;
  reg [31:0] _T_6011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11591;
  reg [31:0] _T_6012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11592;
  reg [31:0] _T_6012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11593;
  reg [31:0] _T_6013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11594;
  reg [31:0] _T_6013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11595;
  reg [31:0] _T_6014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11596;
  reg [31:0] _T_6014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11597;
  reg [31:0] _T_6015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11598;
  reg [31:0] _T_6015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11599;
  reg [31:0] _T_6016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11600;
  reg [31:0] _T_6016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11601;
  reg [31:0] _T_6017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11602;
  reg [31:0] _T_6017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11603;
  reg [31:0] _T_6018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11604;
  reg [31:0] _T_6018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11605;
  reg [31:0] _T_6019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11606;
  reg [31:0] _T_6019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11607;
  reg [31:0] _T_6020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11608;
  reg [31:0] _T_6020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11609;
  reg [31:0] _T_6021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11610;
  reg [31:0] _T_6021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11611;
  reg [31:0] _T_6022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11612;
  reg [31:0] _T_6022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11613;
  reg [31:0] _T_6023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11614;
  reg [31:0] _T_6023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11615;
  reg [31:0] _T_6024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11616;
  reg [31:0] _T_6024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11617;
  reg [31:0] _T_6025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11618;
  reg [31:0] _T_6025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11619;
  reg [31:0] _T_6026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11620;
  reg [31:0] _T_6026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11621;
  reg [31:0] _T_6027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11622;
  reg [31:0] _T_6027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11623;
  reg [31:0] _T_6028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11624;
  reg [31:0] _T_6028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11625;
  reg [31:0] _T_6029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11626;
  reg [31:0] _T_6029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11627;
  reg [31:0] _T_6030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11628;
  reg [31:0] _T_6030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11629;
  reg [31:0] _T_6031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11630;
  reg [31:0] _T_6031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11631;
  reg [31:0] _T_6032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11632;
  reg [31:0] _T_6032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11633;
  reg [31:0] _T_6033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11634;
  reg [31:0] _T_6033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11635;
  reg [31:0] _T_6034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11636;
  reg [31:0] _T_6034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11637;
  reg [31:0] _T_6035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11638;
  reg [31:0] _T_6035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11639;
  reg [31:0] _T_6036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11640;
  reg [31:0] _T_6036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11641;
  reg [31:0] _T_6037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11642;
  reg [31:0] _T_6037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11643;
  reg [31:0] _T_6038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11644;
  reg [31:0] _T_6038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11645;
  reg [31:0] _T_6039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11646;
  reg [31:0] _T_6039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11647;
  reg [31:0] _T_6040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11648;
  reg [31:0] _T_6040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11649;
  reg [31:0] _T_6041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11650;
  reg [31:0] _T_6041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11651;
  reg [31:0] _T_6042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11652;
  reg [31:0] _T_6042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11653;
  reg [31:0] _T_6043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11654;
  reg [31:0] _T_6043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11655;
  reg [31:0] _T_6044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11656;
  reg [31:0] _T_6044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11657;
  reg [31:0] _T_6045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11658;
  reg [31:0] _T_6045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11659;
  reg [31:0] _T_6046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11660;
  reg [31:0] _T_6046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11661;
  reg [31:0] _T_6047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11662;
  reg [31:0] _T_6047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11663;
  reg [31:0] _T_6048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11664;
  reg [31:0] _T_6048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11665;
  reg [31:0] _T_6049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11666;
  reg [31:0] _T_6049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11667;
  reg [31:0] _T_6050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11668;
  reg [31:0] _T_6050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11669;
  reg [31:0] _T_6051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11670;
  reg [31:0] _T_6051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11671;
  reg [31:0] _T_6052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11672;
  reg [31:0] _T_6052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11673;
  reg [31:0] _T_6053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11674;
  reg [31:0] _T_6053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11675;
  reg [31:0] _T_6054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11676;
  reg [31:0] _T_6054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11677;
  reg [31:0] _T_6055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11678;
  reg [31:0] _T_6055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11679;
  reg [31:0] _T_6056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11680;
  reg [31:0] _T_6056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11681;
  reg [31:0] _T_6057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11682;
  reg [31:0] _T_6057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11683;
  reg [31:0] _T_6058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11684;
  reg [31:0] _T_6058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11685;
  reg [31:0] _T_6059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11686;
  reg [31:0] _T_6059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11687;
  reg [31:0] _T_6060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11688;
  reg [31:0] _T_6060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11689;
  reg [31:0] _T_6061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11690;
  reg [31:0] _T_6061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11691;
  reg [31:0] _T_6062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11692;
  reg [31:0] _T_6062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11693;
  reg [31:0] _T_6063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11694;
  reg [31:0] _T_6063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11695;
  reg [31:0] _T_6064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11696;
  reg [31:0] _T_6064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11697;
  reg [31:0] _T_6065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11698;
  reg [31:0] _T_6065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11699;
  reg [31:0] _T_6066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11700;
  reg [31:0] _T_6066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11701;
  reg [31:0] _T_6067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11702;
  reg [31:0] _T_6067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11703;
  reg [31:0] _T_6068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11704;
  reg [31:0] _T_6068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11705;
  reg [31:0] _T_6069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11706;
  reg [31:0] _T_6069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11707;
  reg [31:0] _T_6070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11708;
  reg [31:0] _T_6070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11709;
  reg [31:0] _T_6071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11710;
  reg [31:0] _T_6071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11711;
  reg [31:0] _T_6072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11712;
  reg [31:0] _T_6072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11713;
  reg [31:0] _T_6073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11714;
  reg [31:0] _T_6073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11715;
  reg [31:0] _T_6074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11716;
  reg [31:0] _T_6074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11717;
  reg [31:0] _T_6075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11718;
  reg [31:0] _T_6075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11719;
  reg [31:0] _T_6076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11720;
  reg [31:0] _T_6076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11721;
  reg [31:0] _T_6077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11722;
  reg [31:0] _T_6077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11723;
  reg [31:0] _T_6078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11724;
  reg [31:0] _T_6078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11725;
  reg [31:0] _T_6079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11726;
  reg [31:0] _T_6079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11727;
  reg [31:0] _T_6080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11728;
  reg [31:0] _T_6080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11729;
  reg [31:0] _T_6081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11730;
  reg [31:0] _T_6081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11731;
  reg [31:0] _T_6082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11732;
  reg [31:0] _T_6082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11733;
  reg [31:0] _T_6083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11734;
  reg [31:0] _T_6083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11735;
  reg [31:0] _T_6084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11736;
  reg [31:0] _T_6084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11737;
  reg [31:0] _T_6085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11738;
  reg [31:0] _T_6085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11739;
  reg [31:0] _T_6086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11740;
  reg [31:0] _T_6086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11741;
  reg [31:0] _T_6087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11742;
  reg [31:0] _T_6087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11743;
  reg [31:0] _T_6088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11744;
  reg [31:0] _T_6088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11745;
  reg [31:0] _T_6089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11746;
  reg [31:0] _T_6089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11747;
  reg [31:0] _T_6090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11748;
  reg [31:0] _T_6090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11749;
  reg [31:0] _T_6091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11750;
  reg [31:0] _T_6091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11751;
  reg [31:0] _T_6092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11752;
  reg [31:0] _T_6092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11753;
  reg [31:0] _T_6093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11754;
  reg [31:0] _T_6093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11755;
  reg [31:0] _T_6094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11756;
  reg [31:0] _T_6094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11757;
  reg [31:0] _T_6095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11758;
  reg [31:0] _T_6095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11759;
  reg [31:0] _T_6096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11760;
  reg [31:0] _T_6096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11761;
  reg [31:0] _T_6097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11762;
  reg [31:0] _T_6097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11763;
  reg [31:0] _T_6098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11764;
  reg [31:0] _T_6098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11765;
  reg [31:0] _T_6099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11766;
  reg [31:0] _T_6099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11767;
  reg [31:0] _T_6100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11768;
  reg [31:0] _T_6100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11769;
  reg [31:0] _T_6101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11770;
  reg [31:0] _T_6101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11771;
  reg [31:0] _T_6102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11772;
  reg [31:0] _T_6102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11773;
  reg [31:0] _T_6103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11774;
  reg [31:0] _T_6103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11775;
  reg [31:0] _T_6104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11776;
  reg [31:0] _T_6104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11777;
  reg [31:0] _T_6107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11778;
  reg [31:0] _T_6107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11779;
  reg [31:0] _T_6108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11780;
  reg [31:0] _T_6108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11781;
  reg [31:0] _T_6109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11782;
  reg [31:0] _T_6109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11783;
  reg [31:0] _T_6110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11784;
  reg [31:0] _T_6110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11785;
  reg [31:0] _T_6111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11786;
  reg [31:0] _T_6111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11787;
  reg [31:0] _T_6112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11788;
  reg [31:0] _T_6112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11789;
  reg [31:0] _T_6113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11790;
  reg [31:0] _T_6113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11791;
  reg [31:0] _T_6114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11792;
  reg [31:0] _T_6114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11793;
  reg [31:0] _T_6115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11794;
  reg [31:0] _T_6115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11795;
  reg [31:0] _T_6116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11796;
  reg [31:0] _T_6116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11797;
  reg [31:0] _T_6117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11798;
  reg [31:0] _T_6117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11799;
  reg [31:0] _T_6118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11800;
  reg [31:0] _T_6118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11801;
  reg [31:0] _T_6119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11802;
  reg [31:0] _T_6119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11803;
  reg [31:0] _T_6120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11804;
  reg [31:0] _T_6120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11805;
  reg [31:0] _T_6121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11806;
  reg [31:0] _T_6121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11807;
  reg [31:0] _T_6122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11808;
  reg [31:0] _T_6122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11809;
  reg [31:0] _T_6123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11810;
  reg [31:0] _T_6123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11811;
  reg [31:0] _T_6124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11812;
  reg [31:0] _T_6124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11813;
  reg [31:0] _T_6125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11814;
  reg [31:0] _T_6125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11815;
  reg [31:0] _T_6126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11816;
  reg [31:0] _T_6126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11817;
  reg [31:0] _T_6127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11818;
  reg [31:0] _T_6127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11819;
  reg [31:0] _T_6128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11820;
  reg [31:0] _T_6128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11821;
  reg [31:0] _T_6129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11822;
  reg [31:0] _T_6129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11823;
  reg [31:0] _T_6130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11824;
  reg [31:0] _T_6130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11825;
  reg [31:0] _T_6131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11826;
  reg [31:0] _T_6131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11827;
  reg [31:0] _T_6132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11828;
  reg [31:0] _T_6132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11829;
  reg [31:0] _T_6133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11830;
  reg [31:0] _T_6133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11831;
  reg [31:0] _T_6134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11832;
  reg [31:0] _T_6134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11833;
  reg [31:0] _T_6135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11834;
  reg [31:0] _T_6135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11835;
  reg [31:0] _T_6136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11836;
  reg [31:0] _T_6136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11837;
  reg [31:0] _T_6137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11838;
  reg [31:0] _T_6137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11839;
  reg [31:0] _T_6138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11840;
  reg [31:0] _T_6138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11841;
  reg [31:0] _T_6139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11842;
  reg [31:0] _T_6139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11843;
  reg [31:0] _T_6140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11844;
  reg [31:0] _T_6140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11845;
  reg [31:0] _T_6141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11846;
  reg [31:0] _T_6141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11847;
  reg [31:0] _T_6142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11848;
  reg [31:0] _T_6142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11849;
  reg [31:0] _T_6143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11850;
  reg [31:0] _T_6143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11851;
  reg [31:0] _T_6144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11852;
  reg [31:0] _T_6144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11853;
  reg [31:0] _T_6145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11854;
  reg [31:0] _T_6145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11855;
  reg [31:0] _T_6146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11856;
  reg [31:0] _T_6146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11857;
  reg [31:0] _T_6147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11858;
  reg [31:0] _T_6147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11859;
  reg [31:0] _T_6148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11860;
  reg [31:0] _T_6148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11861;
  reg [31:0] _T_6149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11862;
  reg [31:0] _T_6149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11863;
  reg [31:0] _T_6150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11864;
  reg [31:0] _T_6150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11865;
  reg [31:0] _T_6151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11866;
  reg [31:0] _T_6151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11867;
  reg [31:0] _T_6152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11868;
  reg [31:0] _T_6152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11869;
  reg [31:0] _T_6153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11870;
  reg [31:0] _T_6153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11871;
  reg [31:0] _T_6154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11872;
  reg [31:0] _T_6154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11873;
  reg [31:0] _T_6155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11874;
  reg [31:0] _T_6155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11875;
  reg [31:0] _T_6156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11876;
  reg [31:0] _T_6156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11877;
  reg [31:0] _T_6157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11878;
  reg [31:0] _T_6157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11879;
  reg [31:0] _T_6158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11880;
  reg [31:0] _T_6158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11881;
  reg [31:0] _T_6159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11882;
  reg [31:0] _T_6159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11883;
  reg [31:0] _T_6160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11884;
  reg [31:0] _T_6160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11885;
  reg [31:0] _T_6161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11886;
  reg [31:0] _T_6161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11887;
  reg [31:0] _T_6162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11888;
  reg [31:0] _T_6162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11889;
  reg [31:0] _T_6163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11890;
  reg [31:0] _T_6163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11891;
  reg [31:0] _T_6164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11892;
  reg [31:0] _T_6164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11893;
  reg [31:0] _T_6165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11894;
  reg [31:0] _T_6165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11895;
  reg [31:0] _T_6166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11896;
  reg [31:0] _T_6166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11897;
  reg [31:0] _T_6167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11898;
  reg [31:0] _T_6167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11899;
  reg [31:0] _T_6168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11900;
  reg [31:0] _T_6168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11901;
  reg [31:0] _T_6169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11902;
  reg [31:0] _T_6169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11903;
  reg [31:0] _T_6170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11904;
  reg [31:0] _T_6170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11905;
  wire [31:0] _GEN_19842 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19843 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_19842); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19844 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_19843); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19845 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_19844); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19846 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_19845); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19847 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_19846); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19848 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_19847); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19849 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_19848); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19850 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_19849); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19851 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_19850); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19852 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_19851); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19853 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_19852); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19854 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_19853); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19855 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_19854); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19856 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_19855); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19857 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_19856); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19858 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_19857); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19859 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_19858); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19860 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_19859); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19861 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_19860); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19862 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_19861); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19863 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_19862); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19864 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_19863); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19865 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_19864); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19866 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_19865); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19867 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_19866); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19868 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_19867); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19869 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_19868); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19870 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_19869); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19871 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_19870); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19872 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_19871); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19873 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_19872); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19874 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_19873); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19875 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_19874); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19876 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_19875); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19877 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_19876); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19878 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_19877); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19879 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_19878); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19880 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_19879); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19881 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_19880); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19882 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_19881); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19883 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_19882); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19884 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_19883); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19885 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19884); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19886 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_19885); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19887 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_19886); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19888 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_19887); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19889 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_19888); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19890 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_19889); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19891 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_19890); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19892 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_19891); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19893 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_19892); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19894 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_19893); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19895 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_19894); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19896 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_19895); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19897 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_19896); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19898 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_19897); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19899 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_19898); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19900 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_19899); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19901 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_19900); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19902 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_19901); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19903 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_19902); // @[FFT.scala 34:12]
  wire [31:0] _GEN_19906 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19907 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_19906); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19908 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_19907); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19909 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_19908); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19910 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_19909); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19911 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_19910); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19912 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_19911); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19913 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_19912); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19914 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_19913); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19915 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_19914); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19916 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_19915); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19917 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19916); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19918 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_19917); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19919 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_19918); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19920 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_19919); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19921 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_19920); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19922 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_19921); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19923 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_19922); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19924 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_19923); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19925 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_19924); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19926 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_19925); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19927 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_19926); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19928 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_19927); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19929 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_19928); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19930 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_19929); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19931 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_19930); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19932 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_19931); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19933 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_19932); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19934 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_19933); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19935 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_19934); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19936 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_19935); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19937 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_19936); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19938 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_19937); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19939 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_19938); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19940 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_19939); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19941 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_19940); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19942 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_19941); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19943 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_19942); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19944 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_19943); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19945 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_19944); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19946 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_19945); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19947 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_19946); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19948 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_19947); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19949 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_19948); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19950 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_19949); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19951 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_19950); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19952 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_19951); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19953 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_19952); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19954 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_19953); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19955 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_19954); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19956 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_19955); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19957 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_19956); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19958 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_19957); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19959 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_19958); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19960 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_19959); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19961 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_19960); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19962 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_19961); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19963 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_19962); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19964 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_19963); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19965 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_19964); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19966 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_19965); // @[FFT.scala 35:12]
  wire [31:0] _GEN_19967 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_19966); // @[FFT.scala 35:12]
  reg [31:0] _T_6176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11906;
  reg [31:0] _T_6176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11907;
  reg [31:0] _T_6177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11908;
  reg [31:0] _T_6177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11909;
  reg [31:0] _T_6178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11910;
  reg [31:0] _T_6178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11911;
  reg [31:0] _T_6179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11912;
  reg [31:0] _T_6179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11913;
  reg [31:0] _T_6180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11914;
  reg [31:0] _T_6180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11915;
  reg [31:0] _T_6181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11916;
  reg [31:0] _T_6181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11917;
  reg [31:0] _T_6182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11918;
  reg [31:0] _T_6182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11919;
  reg [31:0] _T_6183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11920;
  reg [31:0] _T_6183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11921;
  reg [31:0] _T_6184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11922;
  reg [31:0] _T_6184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11923;
  reg [31:0] _T_6185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11924;
  reg [31:0] _T_6185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11925;
  reg [31:0] _T_6186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11926;
  reg [31:0] _T_6186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11927;
  reg [31:0] _T_6187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11928;
  reg [31:0] _T_6187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11929;
  reg [31:0] _T_6188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11930;
  reg [31:0] _T_6188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11931;
  reg [31:0] _T_6189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11932;
  reg [31:0] _T_6189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11933;
  reg [31:0] _T_6190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11934;
  reg [31:0] _T_6190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11935;
  reg [31:0] _T_6191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11936;
  reg [31:0] _T_6191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11937;
  reg [31:0] _T_6192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11938;
  reg [31:0] _T_6192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11939;
  reg [31:0] _T_6193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11940;
  reg [31:0] _T_6193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11941;
  reg [31:0] _T_6194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11942;
  reg [31:0] _T_6194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11943;
  reg [31:0] _T_6195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11944;
  reg [31:0] _T_6195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11945;
  reg [31:0] _T_6196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11946;
  reg [31:0] _T_6196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11947;
  reg [31:0] _T_6197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11948;
  reg [31:0] _T_6197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11949;
  reg [31:0] _T_6198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11950;
  reg [31:0] _T_6198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11951;
  reg [31:0] _T_6199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11952;
  reg [31:0] _T_6199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11953;
  reg [31:0] _T_6200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11954;
  reg [31:0] _T_6200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11955;
  reg [31:0] _T_6201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11956;
  reg [31:0] _T_6201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11957;
  reg [31:0] _T_6202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11958;
  reg [31:0] _T_6202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11959;
  reg [31:0] _T_6203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11960;
  reg [31:0] _T_6203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11961;
  reg [31:0] _T_6204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11962;
  reg [31:0] _T_6204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11963;
  reg [31:0] _T_6205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11964;
  reg [31:0] _T_6205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11965;
  reg [31:0] _T_6206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11966;
  reg [31:0] _T_6206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11967;
  reg [31:0] _T_6207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11968;
  reg [31:0] _T_6207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11969;
  reg [31:0] _T_6208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11970;
  reg [31:0] _T_6208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11971;
  reg [31:0] _T_6209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11972;
  reg [31:0] _T_6209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11973;
  reg [31:0] _T_6210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11974;
  reg [31:0] _T_6210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11975;
  reg [31:0] _T_6211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11976;
  reg [31:0] _T_6211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11977;
  reg [31:0] _T_6212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11978;
  reg [31:0] _T_6212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11979;
  reg [31:0] _T_6213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11980;
  reg [31:0] _T_6213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11981;
  reg [31:0] _T_6214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11982;
  reg [31:0] _T_6214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11983;
  reg [31:0] _T_6215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11984;
  reg [31:0] _T_6215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11985;
  reg [31:0] _T_6216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11986;
  reg [31:0] _T_6216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11987;
  reg [31:0] _T_6217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11988;
  reg [31:0] _T_6217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11989;
  reg [31:0] _T_6218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11990;
  reg [31:0] _T_6218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11991;
  reg [31:0] _T_6219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11992;
  reg [31:0] _T_6219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11993;
  reg [31:0] _T_6220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11994;
  reg [31:0] _T_6220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11995;
  reg [31:0] _T_6221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11996;
  reg [31:0] _T_6221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11997;
  reg [31:0] _T_6222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11998;
  reg [31:0] _T_6222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11999;
  reg [31:0] _T_6223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12000;
  reg [31:0] _T_6223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12001;
  reg [31:0] _T_6224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12002;
  reg [31:0] _T_6224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12003;
  reg [31:0] _T_6225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12004;
  reg [31:0] _T_6225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12005;
  reg [31:0] _T_6226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12006;
  reg [31:0] _T_6226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12007;
  reg [31:0] _T_6227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12008;
  reg [31:0] _T_6227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12009;
  reg [31:0] _T_6228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12010;
  reg [31:0] _T_6228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12011;
  reg [31:0] _T_6229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12012;
  reg [31:0] _T_6229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12013;
  reg [31:0] _T_6230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12014;
  reg [31:0] _T_6230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12015;
  reg [31:0] _T_6231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12016;
  reg [31:0] _T_6231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12017;
  reg [31:0] _T_6232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12018;
  reg [31:0] _T_6232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12019;
  reg [31:0] _T_6233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12020;
  reg [31:0] _T_6233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12021;
  reg [31:0] _T_6234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12022;
  reg [31:0] _T_6234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12023;
  reg [31:0] _T_6235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12024;
  reg [31:0] _T_6235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12025;
  reg [31:0] _T_6236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12026;
  reg [31:0] _T_6236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12027;
  reg [31:0] _T_6237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12028;
  reg [31:0] _T_6237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12029;
  reg [31:0] _T_6238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12030;
  reg [31:0] _T_6238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12031;
  reg [31:0] _T_6239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12032;
  reg [31:0] _T_6239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12033;
  reg [31:0] _T_6242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12034;
  reg [31:0] _T_6242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12035;
  reg [31:0] _T_6243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12036;
  reg [31:0] _T_6243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12037;
  reg [31:0] _T_6244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12038;
  reg [31:0] _T_6244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12039;
  reg [31:0] _T_6245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12040;
  reg [31:0] _T_6245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12041;
  reg [31:0] _T_6246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12042;
  reg [31:0] _T_6246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12043;
  reg [31:0] _T_6247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12044;
  reg [31:0] _T_6247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12045;
  reg [31:0] _T_6248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12046;
  reg [31:0] _T_6248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12047;
  reg [31:0] _T_6249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12048;
  reg [31:0] _T_6249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12049;
  reg [31:0] _T_6250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12050;
  reg [31:0] _T_6250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12051;
  reg [31:0] _T_6251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12052;
  reg [31:0] _T_6251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12053;
  reg [31:0] _T_6252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12054;
  reg [31:0] _T_6252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12055;
  reg [31:0] _T_6253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12056;
  reg [31:0] _T_6253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12057;
  reg [31:0] _T_6254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12058;
  reg [31:0] _T_6254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12059;
  reg [31:0] _T_6255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12060;
  reg [31:0] _T_6255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12061;
  reg [31:0] _T_6256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12062;
  reg [31:0] _T_6256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12063;
  reg [31:0] _T_6257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12064;
  reg [31:0] _T_6257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12065;
  reg [31:0] _T_6258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12066;
  reg [31:0] _T_6258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12067;
  reg [31:0] _T_6259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12068;
  reg [31:0] _T_6259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12069;
  reg [31:0] _T_6260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12070;
  reg [31:0] _T_6260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12071;
  reg [31:0] _T_6261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12072;
  reg [31:0] _T_6261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12073;
  reg [31:0] _T_6262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12074;
  reg [31:0] _T_6262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12075;
  reg [31:0] _T_6263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12076;
  reg [31:0] _T_6263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12077;
  reg [31:0] _T_6264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12078;
  reg [31:0] _T_6264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12079;
  reg [31:0] _T_6265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12080;
  reg [31:0] _T_6265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12081;
  reg [31:0] _T_6266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12082;
  reg [31:0] _T_6266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12083;
  reg [31:0] _T_6267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12084;
  reg [31:0] _T_6267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12085;
  reg [31:0] _T_6268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12086;
  reg [31:0] _T_6268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12087;
  reg [31:0] _T_6269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12088;
  reg [31:0] _T_6269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12089;
  reg [31:0] _T_6270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12090;
  reg [31:0] _T_6270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12091;
  reg [31:0] _T_6271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12092;
  reg [31:0] _T_6271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12093;
  reg [31:0] _T_6272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12094;
  reg [31:0] _T_6272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12095;
  reg [31:0] _T_6273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12096;
  reg [31:0] _T_6273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12097;
  wire [31:0] _GEN_20162 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20163 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_20162); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20164 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_20163); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20165 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_20164); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20166 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_20165); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20167 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_20166); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20168 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_20167); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20169 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_20168); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20170 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_20169); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20171 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_20170); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20172 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_20171); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20173 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_20172); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20174 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_20173); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20175 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_20174); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20176 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_20175); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20177 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_20176); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20178 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_20177); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20179 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_20178); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20180 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_20179); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20181 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_20180); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20182 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_20181); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20183 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20182); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20184 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_20183); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20185 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_20184); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20186 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_20185); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20187 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_20186); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20188 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_20187); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20189 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_20188); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20190 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_20189); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20191 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_20190); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20194 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20195 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_20194); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20196 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_20195); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20197 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_20196); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20198 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_20197); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20199 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20198); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20200 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_20199); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20201 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_20200); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20202 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_20201); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20203 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_20202); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20204 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_20203); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20205 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_20204); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20206 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_20205); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20207 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_20206); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20208 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_20207); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20209 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_20208); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20210 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_20209); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20211 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_20210); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20212 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_20211); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20213 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_20212); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20214 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_20213); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20215 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_20214); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20216 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_20215); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20217 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_20216); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20218 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_20217); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20219 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20218); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20220 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_20219); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20221 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_20220); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20222 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_20221); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20223 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_20222); // @[FFT.scala 35:12]
  reg [31:0] _T_6279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12098;
  reg [31:0] _T_6279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12099;
  reg [31:0] _T_6280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12100;
  reg [31:0] _T_6280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12101;
  reg [31:0] _T_6281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12102;
  reg [31:0] _T_6281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12103;
  reg [31:0] _T_6282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12104;
  reg [31:0] _T_6282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12105;
  reg [31:0] _T_6283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12106;
  reg [31:0] _T_6283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12107;
  reg [31:0] _T_6284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12108;
  reg [31:0] _T_6284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12109;
  reg [31:0] _T_6285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12110;
  reg [31:0] _T_6285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12111;
  reg [31:0] _T_6286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12112;
  reg [31:0] _T_6286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12113;
  reg [31:0] _T_6287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12114;
  reg [31:0] _T_6287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12115;
  reg [31:0] _T_6288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12116;
  reg [31:0] _T_6288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12117;
  reg [31:0] _T_6289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12118;
  reg [31:0] _T_6289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12119;
  reg [31:0] _T_6290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12120;
  reg [31:0] _T_6290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12121;
  reg [31:0] _T_6291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12122;
  reg [31:0] _T_6291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12123;
  reg [31:0] _T_6292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12124;
  reg [31:0] _T_6292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12125;
  reg [31:0] _T_6293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12126;
  reg [31:0] _T_6293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12127;
  reg [31:0] _T_6294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12128;
  reg [31:0] _T_6294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12129;
  reg [31:0] _T_6295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12130;
  reg [31:0] _T_6295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12131;
  reg [31:0] _T_6296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12132;
  reg [31:0] _T_6296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12133;
  reg [31:0] _T_6297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12134;
  reg [31:0] _T_6297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12135;
  reg [31:0] _T_6298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12136;
  reg [31:0] _T_6298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12137;
  reg [31:0] _T_6299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12138;
  reg [31:0] _T_6299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12139;
  reg [31:0] _T_6300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12140;
  reg [31:0] _T_6300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12141;
  reg [31:0] _T_6301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12142;
  reg [31:0] _T_6301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12143;
  reg [31:0] _T_6302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12144;
  reg [31:0] _T_6302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12145;
  reg [31:0] _T_6303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12146;
  reg [31:0] _T_6303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12147;
  reg [31:0] _T_6304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12148;
  reg [31:0] _T_6304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12149;
  reg [31:0] _T_6305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12150;
  reg [31:0] _T_6305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12151;
  reg [31:0] _T_6306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12152;
  reg [31:0] _T_6306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12153;
  reg [31:0] _T_6307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12154;
  reg [31:0] _T_6307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12155;
  reg [31:0] _T_6308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12156;
  reg [31:0] _T_6308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12157;
  reg [31:0] _T_6309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12158;
  reg [31:0] _T_6309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12159;
  reg [31:0] _T_6310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12160;
  reg [31:0] _T_6310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12161;
  reg [31:0] _T_6313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12162;
  reg [31:0] _T_6313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12163;
  reg [31:0] _T_6314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12164;
  reg [31:0] _T_6314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12165;
  reg [31:0] _T_6315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12166;
  reg [31:0] _T_6315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12167;
  reg [31:0] _T_6316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12168;
  reg [31:0] _T_6316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12169;
  reg [31:0] _T_6317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12170;
  reg [31:0] _T_6317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12171;
  reg [31:0] _T_6318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12172;
  reg [31:0] _T_6318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12173;
  reg [31:0] _T_6319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12174;
  reg [31:0] _T_6319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12175;
  reg [31:0] _T_6320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12176;
  reg [31:0] _T_6320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12177;
  reg [31:0] _T_6321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12178;
  reg [31:0] _T_6321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12179;
  reg [31:0] _T_6322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12180;
  reg [31:0] _T_6322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12181;
  reg [31:0] _T_6323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12182;
  reg [31:0] _T_6323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12183;
  reg [31:0] _T_6324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12184;
  reg [31:0] _T_6324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12185;
  reg [31:0] _T_6325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12186;
  reg [31:0] _T_6325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12187;
  reg [31:0] _T_6326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12188;
  reg [31:0] _T_6326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12189;
  reg [31:0] _T_6327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12190;
  reg [31:0] _T_6327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12191;
  reg [31:0] _T_6328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12192;
  reg [31:0] _T_6328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12193;
  wire [31:0] _GEN_20322 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20323 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_20322); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20324 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_20323); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20325 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_20324); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20326 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_20325); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20327 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_20326); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20328 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_20327); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20329 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_20328); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20330 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_20329); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20331 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_20330); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20332 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20331); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20333 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_20332); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20334 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_20333); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20335 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_20334); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20338 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20339 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_20338); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20340 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20339); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20341 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_20340); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20342 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_20341); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20343 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_20342); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20344 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_20343); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20345 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_20344); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20346 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_20345); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20347 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_20346); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20348 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_20347); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20349 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_20348); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20350 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_20349); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20351 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_20350); // @[FFT.scala 35:12]
  reg [31:0] _T_6334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12194;
  reg [31:0] _T_6334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12195;
  reg [31:0] _T_6335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12196;
  reg [31:0] _T_6335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12197;
  reg [31:0] _T_6336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12198;
  reg [31:0] _T_6336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12199;
  reg [31:0] _T_6337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12200;
  reg [31:0] _T_6337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12201;
  reg [31:0] _T_6338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12202;
  reg [31:0] _T_6338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12203;
  reg [31:0] _T_6339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12204;
  reg [31:0] _T_6339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12205;
  reg [31:0] _T_6340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12206;
  reg [31:0] _T_6340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12207;
  reg [31:0] _T_6341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12208;
  reg [31:0] _T_6341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12209;
  reg [31:0] _T_6342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12210;
  reg [31:0] _T_6342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12211;
  reg [31:0] _T_6343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12212;
  reg [31:0] _T_6343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12213;
  reg [31:0] _T_6344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12214;
  reg [31:0] _T_6344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12215;
  reg [31:0] _T_6345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12216;
  reg [31:0] _T_6345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12217;
  reg [31:0] _T_6346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12218;
  reg [31:0] _T_6346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12219;
  reg [31:0] _T_6347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12220;
  reg [31:0] _T_6347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12221;
  reg [31:0] _T_6348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12222;
  reg [31:0] _T_6348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12223;
  reg [31:0] _T_6349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12224;
  reg [31:0] _T_6349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12225;
  reg [31:0] _T_6352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12226;
  reg [31:0] _T_6352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12227;
  reg [31:0] _T_6353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12228;
  reg [31:0] _T_6353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12229;
  reg [31:0] _T_6354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12230;
  reg [31:0] _T_6354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12231;
  reg [31:0] _T_6355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12232;
  reg [31:0] _T_6355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12233;
  reg [31:0] _T_6356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12234;
  reg [31:0] _T_6356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12235;
  reg [31:0] _T_6357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12236;
  reg [31:0] _T_6357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12237;
  reg [31:0] _T_6358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12238;
  reg [31:0] _T_6358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12239;
  reg [31:0] _T_6359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12240;
  reg [31:0] _T_6359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12241;
  wire [31:0] _GEN_20402 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20403 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_20402); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20404 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_20403); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20405 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_20404); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20406 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_20405); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20407 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_20406); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20410 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20411 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_20410); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20412 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_20411); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20413 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_20412); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20414 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_20413); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20415 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_20414); // @[FFT.scala 35:12]
  reg [31:0] _T_6365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12242;
  reg [31:0] _T_6365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12243;
  reg [31:0] _T_6366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12244;
  reg [31:0] _T_6366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12245;
  reg [31:0] _T_6367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12246;
  reg [31:0] _T_6367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12247;
  reg [31:0] _T_6368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12248;
  reg [31:0] _T_6368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12249;
  reg [31:0] _T_6369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12250;
  reg [31:0] _T_6369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12251;
  reg [31:0] _T_6370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12252;
  reg [31:0] _T_6370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12253;
  reg [31:0] _T_6371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12254;
  reg [31:0] _T_6371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12255;
  reg [31:0] _T_6372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12256;
  reg [31:0] _T_6372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12257;
  reg [31:0] _T_6375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12258;
  reg [31:0] _T_6375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12259;
  reg [31:0] _T_6376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12260;
  reg [31:0] _T_6376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12261;
  reg [31:0] _T_6377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12262;
  reg [31:0] _T_6377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12263;
  reg [31:0] _T_6378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12264;
  reg [31:0] _T_6378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12265;
  wire [31:0] _GEN_20442 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20443 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_20442); // @[FFT.scala 34:12]
  wire [31:0] _GEN_20446 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  wire [31:0] _GEN_20447 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_20446); // @[FFT.scala 35:12]
  reg [31:0] _T_6384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12266;
  reg [31:0] _T_6384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12267;
  reg [31:0] _T_6385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12268;
  reg [31:0] _T_6385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12269;
  reg [31:0] _T_6386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12270;
  reg [31:0] _T_6386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12271;
  reg [31:0] _T_6387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12272;
  reg [31:0] _T_6387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12273;
  reg [31:0] _T_6390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12274;
  reg [31:0] _T_6390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12275;
  reg [31:0] _T_6391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12276;
  reg [31:0] _T_6391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12277;
  reg [31:0] _T_6397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12278;
  reg [31:0] _T_6397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12279;
  reg [31:0] _T_6398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12280;
  reg [31:0] _T_6398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12281;
  reg [31:0] _T_6401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12282;
  reg [31:0] _T_6401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12283;
  reg [31:0] out1D1_re; // @[FFT.scala 81:23]
  reg [31:0] _RAND_12284;
  reg [31:0] out1D1_im; // @[FFT.scala 81:23]
  reg [31:0] _RAND_12285;
  reg [31:0] _T_6402_re; // @[FFT.scala 85:22]
  reg [31:0] _RAND_12286;
  reg [31:0] _T_6402_im; // @[FFT.scala 85:22]
  reg [31:0] _RAND_12287;
  reg [31:0] _T_6403_re; // @[FFT.scala 86:22]
  reg [31:0] _RAND_12288;
  reg [31:0] _T_6403_im; // @[FFT.scala 86:22]
  reg [31:0] _RAND_12289;
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  Butterfly Butterfly_8 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_8_io_in1_re),
    .io_in1_im(Butterfly_8_io_in1_im),
    .io_in2_re(Butterfly_8_io_in2_re),
    .io_in2_im(Butterfly_8_io_in2_im),
    .io_wn_re(Butterfly_8_io_wn_re),
    .io_wn_im(Butterfly_8_io_wn_im),
    .io_out1_re(Butterfly_8_io_out1_re),
    .io_out1_im(Butterfly_8_io_out1_im),
    .io_out2_re(Butterfly_8_io_out2_re),
    .io_out2_im(Butterfly_8_io_out2_im)
  );
  Switch Switch_8 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_8_io_in1_re),
    .io_in1_im(Switch_8_io_in1_im),
    .io_in2_re(Switch_8_io_in2_re),
    .io_in2_im(Switch_8_io_in2_im),
    .io_sel(Switch_8_io_sel),
    .io_out1_re(Switch_8_io_out1_re),
    .io_out1_im(Switch_8_io_out1_im),
    .io_out2_re(Switch_8_io_out2_re),
    .io_out2_im(Switch_8_io_out2_im)
  );
  Butterfly Butterfly_9 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_9_io_in1_re),
    .io_in1_im(Butterfly_9_io_in1_im),
    .io_in2_re(Butterfly_9_io_in2_re),
    .io_in2_im(Butterfly_9_io_in2_im),
    .io_wn_re(Butterfly_9_io_wn_re),
    .io_wn_im(Butterfly_9_io_wn_im),
    .io_out1_re(Butterfly_9_io_out1_re),
    .io_out1_im(Butterfly_9_io_out1_im),
    .io_out2_re(Butterfly_9_io_out2_re),
    .io_out2_im(Butterfly_9_io_out2_im)
  );
  Switch Switch_9 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_9_io_in1_re),
    .io_in1_im(Switch_9_io_in1_im),
    .io_in2_re(Switch_9_io_in2_re),
    .io_in2_im(Switch_9_io_in2_im),
    .io_sel(Switch_9_io_sel),
    .io_out1_re(Switch_9_io_out1_re),
    .io_out1_im(Switch_9_io_out1_im),
    .io_out2_re(Switch_9_io_out2_re),
    .io_out2_im(Switch_9_io_out2_im)
  );
  Butterfly Butterfly_10 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_10_io_in1_re),
    .io_in1_im(Butterfly_10_io_in1_im),
    .io_in2_re(Butterfly_10_io_in2_re),
    .io_in2_im(Butterfly_10_io_in2_im),
    .io_wn_re(Butterfly_10_io_wn_re),
    .io_wn_im(Butterfly_10_io_wn_im),
    .io_out1_re(Butterfly_10_io_out1_re),
    .io_out1_im(Butterfly_10_io_out1_im),
    .io_out2_re(Butterfly_10_io_out2_re),
    .io_out2_im(Butterfly_10_io_out2_im)
  );
  Switch Switch_10 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_10_io_in1_re),
    .io_in1_im(Switch_10_io_in1_im),
    .io_in2_re(Switch_10_io_in2_re),
    .io_in2_im(Switch_10_io_in2_im),
    .io_sel(Switch_10_io_sel),
    .io_out1_re(Switch_10_io_out1_re),
    .io_out1_im(Switch_10_io_out1_im),
    .io_out2_re(Switch_10_io_out2_re),
    .io_out2_im(Switch_10_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign io_dOut1_re = _T_6402_re; // @[FFT.scala 85:12]
  assign io_dOut1_im = _T_6402_im; // @[FFT.scala 85:12]
  assign io_dOut2_re = _T_6403_re; // @[FFT.scala 86:12]
  assign io_dOut2_im = _T_6403_im; // @[FFT.scala 86:12]
  assign io_dout_valid = cntD1 == 12'hfff; // @[FFT.scala 91:19]
  assign Butterfly_io_in1_re = _T_2236_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_2236_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 11'h7ff == cnt[10:0] ? $signed(-32'sh10000) : $signed(_GEN_2047); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 11'h7ff == cnt[10:0] ? $signed(-32'sh65) : $signed(_GEN_4095); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_3262_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_3262_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[10]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_4291_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_4291_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 10'h3ff == cnt[9:0] ? $signed(-32'sh10000) : $signed(_GEN_11263); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 10'h3ff == cnt[9:0] ? $signed(-32'shc9) : $signed(_GEN_12287); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_4805_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_4805_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[9]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_5322_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_5322_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 9'h1ff == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_15871); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 9'h1ff == cnt[8:0] ? $signed(-32'sh192) : $signed(_GEN_16383); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_5580_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_5580_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[8]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_5841_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_5841_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 8'hff == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_18175); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 8'hff == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_18431); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_5971_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_5971_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[7]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_6104_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_6104_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_19327); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_19455); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_6170_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_6170_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[6]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_6239_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_6239_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_19903); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_19967); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_6273_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_6273_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_6310_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_6310_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_20191); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_20223); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_6328_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_6328_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_6349_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_6349_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_20335); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_20351); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_6359_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_6359_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_8_io_in1_re = _T_6372_re; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in1_im = _T_6372_im; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in2_re = Switch_7_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_in2_im = Switch_7_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_20407); // @[Butterfly.scala 92:16]
  assign Butterfly_8_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_20415); // @[Butterfly.scala 92:16]
  assign Switch_8_io_in1_re = Butterfly_8_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in1_im = Butterfly_8_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in2_re = _T_6378_re; // @[Butterfly.scala 112:17]
  assign Switch_8_io_in2_im = _T_6378_im; // @[Butterfly.scala 112:17]
  assign Switch_8_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_9_io_in1_re = _T_6387_re; // @[Butterfly.scala 90:17]
  assign Butterfly_9_io_in1_im = _T_6387_im; // @[Butterfly.scala 90:17]
  assign Butterfly_9_io_in2_re = Switch_8_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_9_io_in2_im = Switch_8_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_9_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_20443); // @[Butterfly.scala 92:16]
  assign Butterfly_9_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_20447); // @[Butterfly.scala 92:16]
  assign Switch_9_io_in1_re = Butterfly_9_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_9_io_in1_im = Butterfly_9_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_9_io_in2_re = _T_6391_re; // @[Butterfly.scala 112:17]
  assign Switch_9_io_in2_im = _T_6391_im; // @[Butterfly.scala 112:17]
  assign Switch_9_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_10_io_in1_re = _T_6398_re; // @[Butterfly.scala 90:17]
  assign Butterfly_10_io_in1_im = _T_6398_im; // @[Butterfly.scala 90:17]
  assign Butterfly_10_io_in2_re = Switch_9_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_10_io_in2_im = Switch_9_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_10_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_10_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_10_io_in1_re = Butterfly_10_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_10_io_in1_im = Butterfly_10_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_10_io_in2_re = _T_6401_re; // @[Butterfly.scala 112:17]
  assign Switch_10_io_in2_im = _T_6401_im; // @[Butterfly.scala 112:17]
  assign Switch_10_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_10_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_10_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_10_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_10_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntD1 = _RAND_1[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_189_re = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_189_im = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_190_re = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_190_im = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_191_re = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_191_im = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_192_re = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_192_im = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_193_re = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_193_im = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_194_re = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_194_im = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_195_re = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_195_im = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_196_re = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_196_im = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_197_re = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_197_im = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_198_re = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_198_im = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_199_re = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_199_im = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_200_re = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_200_im = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_201_re = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_201_im = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_202_re = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_202_im = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_203_re = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_203_im = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_204_re = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_204_im = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_205_re = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_205_im = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_206_re = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_206_im = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_207_re = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_207_im = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_208_re = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_208_im = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_209_re = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_209_im = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_210_re = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_210_im = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_211_re = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_211_im = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_212_re = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_212_im = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_213_re = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_213_im = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_214_re = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_214_im = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_215_re = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_215_im = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_216_re = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_216_im = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_217_re = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_217_im = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_218_re = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_218_im = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_219_re = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_219_im = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_220_re = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_220_im = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_221_re = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_221_im = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_222_re = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_222_im = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_223_re = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_223_im = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_224_re = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_224_im = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_225_re = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_225_im = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_226_re = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_226_im = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_227_re = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_227_im = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_228_re = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_228_im = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_229_re = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_229_im = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_230_re = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_230_im = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_231_re = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_231_im = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_232_re = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_232_im = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_233_re = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_233_im = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_234_re = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_234_im = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_235_re = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_235_im = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_236_re = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_236_im = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_237_re = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_237_im = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_238_re = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_238_im = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_239_re = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_239_im = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_240_re = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_240_im = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_241_re = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_241_im = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_242_re = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_242_im = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_243_re = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_243_im = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_244_re = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_244_im = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_245_re = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_245_im = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_246_re = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_246_im = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_247_re = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_247_im = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_248_re = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_248_im = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_249_re = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_249_im = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_250_re = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_250_im = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_251_re = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_251_im = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_252_re = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_252_im = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_253_re = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_253_im = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_254_re = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_254_im = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_255_re = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_255_im = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_256_re = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_256_im = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_257_re = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_257_im = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_258_re = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_258_im = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_259_re = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_259_im = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_260_re = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_260_im = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_261_re = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_261_im = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_262_re = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_262_im = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_263_re = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_263_im = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_264_re = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_264_im = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_265_re = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_265_im = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_266_re = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_266_im = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_267_re = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_267_im = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_268_re = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_268_im = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_269_re = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_269_im = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_270_re = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_270_im = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_271_re = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_271_im = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_272_re = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_272_im = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_273_re = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_273_im = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_274_re = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_274_im = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_275_re = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_275_im = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_276_re = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_276_im = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_277_re = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_277_im = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_278_re = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_278_im = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_279_re = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_279_im = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_280_re = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_280_im = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_281_re = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_281_im = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_282_re = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_282_im = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_283_re = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_283_im = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_284_re = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_284_im = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_285_re = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_285_im = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_286_re = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_286_im = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_287_re = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_287_im = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_288_re = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_288_im = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_289_re = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_289_im = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_290_re = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_290_im = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_291_re = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_291_im = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_292_re = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_292_im = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_293_re = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_293_im = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_294_re = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_294_im = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_295_re = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_295_im = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_296_re = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_296_im = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_297_re = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_297_im = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_298_re = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_298_im = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_299_re = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_299_im = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_300_re = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_300_im = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_301_re = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_301_im = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_302_re = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_302_im = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_303_re = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_303_im = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_304_re = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_304_im = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_305_re = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_305_im = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_306_re = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_306_im = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_307_re = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_307_im = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_308_re = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_308_im = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_309_re = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_309_im = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_310_re = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_310_im = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_311_re = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_311_im = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_312_re = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_312_im = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_313_re = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_313_im = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_314_re = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_314_im = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_315_re = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_315_im = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_316_re = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_316_im = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_317_re = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_317_im = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_318_re = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_318_im = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_319_re = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_319_im = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_320_re = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_320_im = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_321_re = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_321_im = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_322_re = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_322_im = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_323_re = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_323_im = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_324_re = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_324_im = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_325_re = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_325_im = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_326_re = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_326_im = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_327_re = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_327_im = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_328_re = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_328_im = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_329_re = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_329_im = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_330_re = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_330_im = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_331_re = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_331_im = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_332_re = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_332_im = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_333_re = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_333_im = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_334_re = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_334_im = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_335_re = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_335_im = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_336_re = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_336_im = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_337_re = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_337_im = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_338_re = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_338_im = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_339_re = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_339_im = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_340_re = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_340_im = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_341_re = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_341_im = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_342_re = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_342_im = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_343_re = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_343_im = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_344_re = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_344_im = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_345_re = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_345_im = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_346_re = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_346_im = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_347_re = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_347_im = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_348_re = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_348_im = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_349_re = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_349_im = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_350_re = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_350_im = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_351_re = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_351_im = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_352_re = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_352_im = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_353_re = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_353_im = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_354_re = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_354_im = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_355_re = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_355_im = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_356_re = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_356_im = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_357_re = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_357_im = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_358_re = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_358_im = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_359_re = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_359_im = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_360_re = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_360_im = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_361_re = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_361_im = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_362_re = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_362_im = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_363_re = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_363_im = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_364_re = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_364_im = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_365_re = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_365_im = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_366_re = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_366_im = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_367_re = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_367_im = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_368_re = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_368_im = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_369_re = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_369_im = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_370_re = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_370_im = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_371_re = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_371_im = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_372_re = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_372_im = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_373_re = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_373_im = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_374_re = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_374_im = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_375_re = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_375_im = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_376_re = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_376_im = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_377_re = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_377_im = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_378_re = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_378_im = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_379_re = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_379_im = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_380_re = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_380_im = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_381_re = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_381_im = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_382_re = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_382_im = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_383_re = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_383_im = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_384_re = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_384_im = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_385_re = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_385_im = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_386_re = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_386_im = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_387_re = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_387_im = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_388_re = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_388_im = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_389_re = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_389_im = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_390_re = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_390_im = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_391_re = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_391_im = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_392_re = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_392_im = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_393_re = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_393_im = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_394_re = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_394_im = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_395_re = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_395_im = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_396_re = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_396_im = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_397_re = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_397_im = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_398_re = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_398_im = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_399_re = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_399_im = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_400_re = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_400_im = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_401_re = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_401_im = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_402_re = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_402_im = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_403_re = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_403_im = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_404_re = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_404_im = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_405_re = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_405_im = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_406_re = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_406_im = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_407_re = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_407_im = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_408_re = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_408_im = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_409_re = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_409_im = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_410_re = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_410_im = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_411_re = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_411_im = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_412_re = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_412_im = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_413_re = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_413_im = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_414_re = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_414_im = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_415_re = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_415_im = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_416_re = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_416_im = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_417_re = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_417_im = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_418_re = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_418_im = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_419_re = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_419_im = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_420_re = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_420_im = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_421_re = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_421_im = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_422_re = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_422_im = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_423_re = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_423_im = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_424_re = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_424_im = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_425_re = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_425_im = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_426_re = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_426_im = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_427_re = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_427_im = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_428_re = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_428_im = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_429_re = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_429_im = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_430_re = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_430_im = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_431_re = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_431_im = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_432_re = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_432_im = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_433_re = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_433_im = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_434_re = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_434_im = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_435_re = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_435_im = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_436_re = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_436_im = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_437_re = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_437_im = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_438_re = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_438_im = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_439_re = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_439_im = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_440_re = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_440_im = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_441_re = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_441_im = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_442_re = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_442_im = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_443_re = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_443_im = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_444_re = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_444_im = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_445_re = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_445_im = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_446_re = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_446_im = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_447_re = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_447_im = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_448_re = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_448_im = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_449_re = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_449_im = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_450_re = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_450_im = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_451_re = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_451_im = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_452_re = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_452_im = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_453_re = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_453_im = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_454_re = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_454_im = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_455_re = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_455_im = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_456_re = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_456_im = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_457_re = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_457_im = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_458_re = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_458_im = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_459_re = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_459_im = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_460_re = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_460_im = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_461_re = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_461_im = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_462_re = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_462_im = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_463_re = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_463_im = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_464_re = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_464_im = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_465_re = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_465_im = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_466_re = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_466_im = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_467_re = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_467_im = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_468_re = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_468_im = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_469_re = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_469_im = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_470_re = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_470_im = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_471_re = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_471_im = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_472_re = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_472_im = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_473_re = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_473_im = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_474_re = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_474_im = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_475_re = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_475_im = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_476_re = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_476_im = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_477_re = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_477_im = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_478_re = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_478_im = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_479_re = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_479_im = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_480_re = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_480_im = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_481_re = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_481_im = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_482_re = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_482_im = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_483_re = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_483_im = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_484_re = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_484_im = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_485_re = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_485_im = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_486_re = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_486_im = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_487_re = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_487_im = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_488_re = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_488_im = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_489_re = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_489_im = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_490_re = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_490_im = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_491_re = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_491_im = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_492_re = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_492_im = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_493_re = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_493_im = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_494_re = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_494_im = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_495_re = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_495_im = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_496_re = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_496_im = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_497_re = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_497_im = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_498_re = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_498_im = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_499_re = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_499_im = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_500_re = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_500_im = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_501_re = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_501_im = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_502_re = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_502_im = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_503_re = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_503_im = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_504_re = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_504_im = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_505_re = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_505_im = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_506_re = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_506_im = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_507_re = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_507_im = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_508_re = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_508_im = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_509_re = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_509_im = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_510_re = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_510_im = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_511_re = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_511_im = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_512_re = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_512_im = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_513_re = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_513_im = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_514_re = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_514_im = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_515_re = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_515_im = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_516_re = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_516_im = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_517_re = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_517_im = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_518_re = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_518_im = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_519_re = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_519_im = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_520_re = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_520_im = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_521_re = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_521_im = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_522_re = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_522_im = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_523_re = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_523_im = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_524_re = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_524_im = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_525_re = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_525_im = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_526_re = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_526_im = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_527_re = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_527_im = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_528_re = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_528_im = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_529_re = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_529_im = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_530_re = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_530_im = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_531_re = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_531_im = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_532_re = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_532_im = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_533_re = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_533_im = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_534_re = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_534_im = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_535_re = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_535_im = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_536_re = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_536_im = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_537_re = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_537_im = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_538_re = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_538_im = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_539_re = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_539_im = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_540_re = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_540_im = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_541_re = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_541_im = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_542_re = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_542_im = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_543_re = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_543_im = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_544_re = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_544_im = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_545_re = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_545_im = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_546_re = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_546_im = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_547_re = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_547_im = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_548_re = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_548_im = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_549_re = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_549_im = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_550_re = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_550_im = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_551_re = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_551_im = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_552_re = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_552_im = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_553_re = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_553_im = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_554_re = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_554_im = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_555_re = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_555_im = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_556_re = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_556_im = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_557_re = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_557_im = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_558_re = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_558_im = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_559_re = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_559_im = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_560_re = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_560_im = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_561_re = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_561_im = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_562_re = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_562_im = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_563_re = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_563_im = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_564_re = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_564_im = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_565_re = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_565_im = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_566_re = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_566_im = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_567_re = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_567_im = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_568_re = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_568_im = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_569_re = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_569_im = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_570_re = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_570_im = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_571_re = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_571_im = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_572_re = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_572_im = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_573_re = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_573_im = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_574_re = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_574_im = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_575_re = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_575_im = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_576_re = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_576_im = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_577_re = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_577_im = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_578_re = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_578_im = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_579_re = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_579_im = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_580_re = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_580_im = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_581_re = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_581_im = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_582_re = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_582_im = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_583_re = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_583_im = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_584_re = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_584_im = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_585_re = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_585_im = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_586_re = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_586_im = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_587_re = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_587_im = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_588_re = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_588_im = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_589_re = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_589_im = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_590_re = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_590_im = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_591_re = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_591_im = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_592_re = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_592_im = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_593_re = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_593_im = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_594_re = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_594_im = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_595_re = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_595_im = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_596_re = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_596_im = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_597_re = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_597_im = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_598_re = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_598_im = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_599_re = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_599_im = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_600_re = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_600_im = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_601_re = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_601_im = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_602_re = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_602_im = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_603_re = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_603_im = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_604_re = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_604_im = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_605_re = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_605_im = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_606_re = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_606_im = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_607_re = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_607_im = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_608_re = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_608_im = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_609_re = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_609_im = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_610_re = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_610_im = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_611_re = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_611_im = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_612_re = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_612_im = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_613_re = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_613_im = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_614_re = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_614_im = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_615_re = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_615_im = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_616_re = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_616_im = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_617_re = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_617_im = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_618_re = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_618_im = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_619_re = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_619_im = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_620_re = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_620_im = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_621_re = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_621_im = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_622_re = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_622_im = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_623_re = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_623_im = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_624_re = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_624_im = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_625_re = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_625_im = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_626_re = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_626_im = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_627_re = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_627_im = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_628_re = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_628_im = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_629_re = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_629_im = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_630_re = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_630_im = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_631_re = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_631_im = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_632_re = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_632_im = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_633_re = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_633_im = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_634_re = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_634_im = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_635_re = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_635_im = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_636_re = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_636_im = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_637_re = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_637_im = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_638_re = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_638_im = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_639_re = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_639_im = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_640_re = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_640_im = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_641_re = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_641_im = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_642_re = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_642_im = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_643_re = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_643_im = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_644_re = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_644_im = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_645_re = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_645_im = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_646_re = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_646_im = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_647_re = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_647_im = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_648_re = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_648_im = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_649_re = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_649_im = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_650_re = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_650_im = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_651_re = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_651_im = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_652_re = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_652_im = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_653_re = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_653_im = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_654_re = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_654_im = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_655_re = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_655_im = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_656_re = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_656_im = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_657_re = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_657_im = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_658_re = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_658_im = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_659_re = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_659_im = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_660_re = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_660_im = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_661_re = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_661_im = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_662_re = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_662_im = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_663_re = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_663_im = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_664_re = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_664_im = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_665_re = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_665_im = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_666_re = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_666_im = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_667_re = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_667_im = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_668_re = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_668_im = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_669_re = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_669_im = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_670_re = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_670_im = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_671_re = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_671_im = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_672_re = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_672_im = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_673_re = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_673_im = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_674_re = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_674_im = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_675_re = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_675_im = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_676_re = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_676_im = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_677_re = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_677_im = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_678_re = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_678_im = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_679_re = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_679_im = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_680_re = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_680_im = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_681_re = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_681_im = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_682_re = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_682_im = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_683_re = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_683_im = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_684_re = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_684_im = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_685_re = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_685_im = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_686_re = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_686_im = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_687_re = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_687_im = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_688_re = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_688_im = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_689_re = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_689_im = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_690_re = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_690_im = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_691_re = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_691_im = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_692_re = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_692_im = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_693_re = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_693_im = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_694_re = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_694_im = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_695_re = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_695_im = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_696_re = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_696_im = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_697_re = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_697_im = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_698_re = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_698_im = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_699_re = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_699_im = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_700_re = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_700_im = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_701_re = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_701_im = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_702_re = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_702_im = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_703_re = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_703_im = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_704_re = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_704_im = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_705_re = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_705_im = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_706_re = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_706_im = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_707_re = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_707_im = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_708_re = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_708_im = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_709_re = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_709_im = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_710_re = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_710_im = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_711_re = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_711_im = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_712_re = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_712_im = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_713_re = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_713_im = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_714_re = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_714_im = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_715_re = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_715_im = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_716_re = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_716_im = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_717_re = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_717_im = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_718_re = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_718_im = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_719_re = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_719_im = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_720_re = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_720_im = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_721_re = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_721_im = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_722_re = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_722_im = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_723_re = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_723_im = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_724_re = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_724_im = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_725_re = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_725_im = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_726_re = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_726_im = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_727_re = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_727_im = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_728_re = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_728_im = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_729_re = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_729_im = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_730_re = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_730_im = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_731_re = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_731_im = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_732_re = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_732_im = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_733_re = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_733_im = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_734_re = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_734_im = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_735_re = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_735_im = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_736_re = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_736_im = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_737_re = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_737_im = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_738_re = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_738_im = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_739_re = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_739_im = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_740_re = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_740_im = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_741_re = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_741_im = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_742_re = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_742_im = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_743_re = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_743_im = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_744_re = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_744_im = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_745_re = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_745_im = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_746_re = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_746_im = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_747_re = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_747_im = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_748_re = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_748_im = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_749_re = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_749_im = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_750_re = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_750_im = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_751_re = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_751_im = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_752_re = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_752_im = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_753_re = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_753_im = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_754_re = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_754_im = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_755_re = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_755_im = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_756_re = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_756_im = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_757_re = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_757_im = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_758_re = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_758_im = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_759_re = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_759_im = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_760_re = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_760_im = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_761_re = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_761_im = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_762_re = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_762_im = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_763_re = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_763_im = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_764_re = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_764_im = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_765_re = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_765_im = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_766_re = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_766_im = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_767_re = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_767_im = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_768_re = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_768_im = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_769_re = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_769_im = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_770_re = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_770_im = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_771_re = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_771_im = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_772_re = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_772_im = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_773_re = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_773_im = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_774_re = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_774_im = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_775_re = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_775_im = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_776_re = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_776_im = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_777_re = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_777_im = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_778_re = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_778_im = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_779_re = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_779_im = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_780_re = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_780_im = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_781_re = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_781_im = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_782_re = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_782_im = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_783_re = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_783_im = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_784_re = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_784_im = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_785_re = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_785_im = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_786_re = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_786_im = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_787_re = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_787_im = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_788_re = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_788_im = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_789_re = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_789_im = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_790_re = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_790_im = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_791_re = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_791_im = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_792_re = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_792_im = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_793_re = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_793_im = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_794_re = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_794_im = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_795_re = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_795_im = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_796_re = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_796_im = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_797_re = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_797_im = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_798_re = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_798_im = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_799_re = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_799_im = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_800_re = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_800_im = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_801_re = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_801_im = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_802_re = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_802_im = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_803_re = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_803_im = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_804_re = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_804_im = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_805_re = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_805_im = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_806_re = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_806_im = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_807_re = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_807_im = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_808_re = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_808_im = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_809_re = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_809_im = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_810_re = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_810_im = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_811_re = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_811_im = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_812_re = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_812_im = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_813_re = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_813_im = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_814_re = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_814_im = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_815_re = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_815_im = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_816_re = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_816_im = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_817_re = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_817_im = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_818_re = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_818_im = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_819_re = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_819_im = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_820_re = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_820_im = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_821_re = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_821_im = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_822_re = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_822_im = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_823_re = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_823_im = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_824_re = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_824_im = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_825_re = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_825_im = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_826_re = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_826_im = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_827_re = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_827_im = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_828_re = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_828_im = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_829_re = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_829_im = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_830_re = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_830_im = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_831_re = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_831_im = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_832_re = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_832_im = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_833_re = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_833_im = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_834_re = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_834_im = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_835_re = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_835_im = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_836_re = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_836_im = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_837_re = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_837_im = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_838_re = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_838_im = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_839_re = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_839_im = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_840_re = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_840_im = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_841_re = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_841_im = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_842_re = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_842_im = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_843_re = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_843_im = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_844_re = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_844_im = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_845_re = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_845_im = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_846_re = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_846_im = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_847_re = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_847_im = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_848_re = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_848_im = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_849_re = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_849_im = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_850_re = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_850_im = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_851_re = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_851_im = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_852_re = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_852_im = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_853_re = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_853_im = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_854_re = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_854_im = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_855_re = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_855_im = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_856_re = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_856_im = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_857_re = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_857_im = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_858_re = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_858_im = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_859_re = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_859_im = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_860_re = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_860_im = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_861_re = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_861_im = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_862_re = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_862_im = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_863_re = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_863_im = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_864_re = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_864_im = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_865_re = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_865_im = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_866_re = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_866_im = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_867_re = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_867_im = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_868_re = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_868_im = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_869_re = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_869_im = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_870_re = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_870_im = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_871_re = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_871_im = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_872_re = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_872_im = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_873_re = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_873_im = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_874_re = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_874_im = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_875_re = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_875_im = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_876_re = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_876_im = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_877_re = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_877_im = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_878_re = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_878_im = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_879_re = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_879_im = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_880_re = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_880_im = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_881_re = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_881_im = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_882_re = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_882_im = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_883_re = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_883_im = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_884_re = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_884_im = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_885_re = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_885_im = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_886_re = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_886_im = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_887_re = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_887_im = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_888_re = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_888_im = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_889_re = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_889_im = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_890_re = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_890_im = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_891_re = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_891_im = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_892_re = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_892_im = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_893_re = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_893_im = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_894_re = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_894_im = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_895_re = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_895_im = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_896_re = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_896_im = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_897_re = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_897_im = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_898_re = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_898_im = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_899_re = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_899_im = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_900_re = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_900_im = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_901_re = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_901_im = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_902_re = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_902_im = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_903_re = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_903_im = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_904_re = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_904_im = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_905_re = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_905_im = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_906_re = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_906_im = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_907_re = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_907_im = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_908_re = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_908_im = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_909_re = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_909_im = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_910_re = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_910_im = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_911_re = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_911_im = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_912_re = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_912_im = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_913_re = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_913_im = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_914_re = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_914_im = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_915_re = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_915_im = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_916_re = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_916_im = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_917_re = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_917_im = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_918_re = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_918_im = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_919_re = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_919_im = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_920_re = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_920_im = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_921_re = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_921_im = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_922_re = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_922_im = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_923_re = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_923_im = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_924_re = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_924_im = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_925_re = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_925_im = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_926_re = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_926_im = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_927_re = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_927_im = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_928_re = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_928_im = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_929_re = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_929_im = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_930_re = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_930_im = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_931_re = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_931_im = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_932_re = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_932_im = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_933_re = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_933_im = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_934_re = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_934_im = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_935_re = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_935_im = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_936_re = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_936_im = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_937_re = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_937_im = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_938_re = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_938_im = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_939_re = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_939_im = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_940_re = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_940_im = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_941_re = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_941_im = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_942_re = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_942_im = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_943_re = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_943_im = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_944_re = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_944_im = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_945_re = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_945_im = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_946_re = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_946_im = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_947_re = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_947_im = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_948_re = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_948_im = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_949_re = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_949_im = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_950_re = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_950_im = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_951_re = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_951_im = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_952_re = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_952_im = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_953_re = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  _T_953_im = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  _T_954_re = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_954_im = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_955_re = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_955_im = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_956_re = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  _T_956_im = _RAND_1537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  _T_957_re = _RAND_1538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_957_im = _RAND_1539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_958_re = _RAND_1540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_958_im = _RAND_1541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_959_re = _RAND_1542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{`RANDOM}};
  _T_959_im = _RAND_1543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{`RANDOM}};
  _T_960_re = _RAND_1544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{`RANDOM}};
  _T_960_im = _RAND_1545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{`RANDOM}};
  _T_961_re = _RAND_1546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{`RANDOM}};
  _T_961_im = _RAND_1547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{`RANDOM}};
  _T_962_re = _RAND_1548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{`RANDOM}};
  _T_962_im = _RAND_1549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{`RANDOM}};
  _T_963_re = _RAND_1550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{`RANDOM}};
  _T_963_im = _RAND_1551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{`RANDOM}};
  _T_964_re = _RAND_1552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{`RANDOM}};
  _T_964_im = _RAND_1553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{`RANDOM}};
  _T_965_re = _RAND_1554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{`RANDOM}};
  _T_965_im = _RAND_1555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{`RANDOM}};
  _T_966_re = _RAND_1556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{`RANDOM}};
  _T_966_im = _RAND_1557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{`RANDOM}};
  _T_967_re = _RAND_1558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{`RANDOM}};
  _T_967_im = _RAND_1559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{`RANDOM}};
  _T_968_re = _RAND_1560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{`RANDOM}};
  _T_968_im = _RAND_1561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{`RANDOM}};
  _T_969_re = _RAND_1562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{`RANDOM}};
  _T_969_im = _RAND_1563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{`RANDOM}};
  _T_970_re = _RAND_1564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{`RANDOM}};
  _T_970_im = _RAND_1565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{`RANDOM}};
  _T_971_re = _RAND_1566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{`RANDOM}};
  _T_971_im = _RAND_1567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{`RANDOM}};
  _T_972_re = _RAND_1568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{`RANDOM}};
  _T_972_im = _RAND_1569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{`RANDOM}};
  _T_973_re = _RAND_1570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{`RANDOM}};
  _T_973_im = _RAND_1571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{`RANDOM}};
  _T_974_re = _RAND_1572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{`RANDOM}};
  _T_974_im = _RAND_1573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{`RANDOM}};
  _T_975_re = _RAND_1574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{`RANDOM}};
  _T_975_im = _RAND_1575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{`RANDOM}};
  _T_976_re = _RAND_1576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{`RANDOM}};
  _T_976_im = _RAND_1577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{`RANDOM}};
  _T_977_re = _RAND_1578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{`RANDOM}};
  _T_977_im = _RAND_1579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{`RANDOM}};
  _T_978_re = _RAND_1580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{`RANDOM}};
  _T_978_im = _RAND_1581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{`RANDOM}};
  _T_979_re = _RAND_1582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{`RANDOM}};
  _T_979_im = _RAND_1583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{`RANDOM}};
  _T_980_re = _RAND_1584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{`RANDOM}};
  _T_980_im = _RAND_1585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{`RANDOM}};
  _T_981_re = _RAND_1586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{`RANDOM}};
  _T_981_im = _RAND_1587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{`RANDOM}};
  _T_982_re = _RAND_1588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{`RANDOM}};
  _T_982_im = _RAND_1589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{`RANDOM}};
  _T_983_re = _RAND_1590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{`RANDOM}};
  _T_983_im = _RAND_1591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{`RANDOM}};
  _T_984_re = _RAND_1592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{`RANDOM}};
  _T_984_im = _RAND_1593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{`RANDOM}};
  _T_985_re = _RAND_1594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{`RANDOM}};
  _T_985_im = _RAND_1595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{`RANDOM}};
  _T_986_re = _RAND_1596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{`RANDOM}};
  _T_986_im = _RAND_1597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{`RANDOM}};
  _T_987_re = _RAND_1598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{`RANDOM}};
  _T_987_im = _RAND_1599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{`RANDOM}};
  _T_988_re = _RAND_1600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{`RANDOM}};
  _T_988_im = _RAND_1601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{`RANDOM}};
  _T_989_re = _RAND_1602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{`RANDOM}};
  _T_989_im = _RAND_1603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{`RANDOM}};
  _T_990_re = _RAND_1604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{`RANDOM}};
  _T_990_im = _RAND_1605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{`RANDOM}};
  _T_991_re = _RAND_1606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{`RANDOM}};
  _T_991_im = _RAND_1607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{`RANDOM}};
  _T_992_re = _RAND_1608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{`RANDOM}};
  _T_992_im = _RAND_1609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{`RANDOM}};
  _T_993_re = _RAND_1610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{`RANDOM}};
  _T_993_im = _RAND_1611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{`RANDOM}};
  _T_994_re = _RAND_1612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{`RANDOM}};
  _T_994_im = _RAND_1613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{`RANDOM}};
  _T_995_re = _RAND_1614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{`RANDOM}};
  _T_995_im = _RAND_1615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{`RANDOM}};
  _T_996_re = _RAND_1616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{`RANDOM}};
  _T_996_im = _RAND_1617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{`RANDOM}};
  _T_997_re = _RAND_1618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{`RANDOM}};
  _T_997_im = _RAND_1619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{`RANDOM}};
  _T_998_re = _RAND_1620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{`RANDOM}};
  _T_998_im = _RAND_1621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{`RANDOM}};
  _T_999_re = _RAND_1622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{`RANDOM}};
  _T_999_im = _RAND_1623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{`RANDOM}};
  _T_1000_re = _RAND_1624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{`RANDOM}};
  _T_1000_im = _RAND_1625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{`RANDOM}};
  _T_1001_re = _RAND_1626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{`RANDOM}};
  _T_1001_im = _RAND_1627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{`RANDOM}};
  _T_1002_re = _RAND_1628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{`RANDOM}};
  _T_1002_im = _RAND_1629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{`RANDOM}};
  _T_1003_re = _RAND_1630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{`RANDOM}};
  _T_1003_im = _RAND_1631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{`RANDOM}};
  _T_1004_re = _RAND_1632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{`RANDOM}};
  _T_1004_im = _RAND_1633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{`RANDOM}};
  _T_1005_re = _RAND_1634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{`RANDOM}};
  _T_1005_im = _RAND_1635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{`RANDOM}};
  _T_1006_re = _RAND_1636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{`RANDOM}};
  _T_1006_im = _RAND_1637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{`RANDOM}};
  _T_1007_re = _RAND_1638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{`RANDOM}};
  _T_1007_im = _RAND_1639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{`RANDOM}};
  _T_1008_re = _RAND_1640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{`RANDOM}};
  _T_1008_im = _RAND_1641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{`RANDOM}};
  _T_1009_re = _RAND_1642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{`RANDOM}};
  _T_1009_im = _RAND_1643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{`RANDOM}};
  _T_1010_re = _RAND_1644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{`RANDOM}};
  _T_1010_im = _RAND_1645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{`RANDOM}};
  _T_1011_re = _RAND_1646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{`RANDOM}};
  _T_1011_im = _RAND_1647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{`RANDOM}};
  _T_1012_re = _RAND_1648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{`RANDOM}};
  _T_1012_im = _RAND_1649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{`RANDOM}};
  _T_1013_re = _RAND_1650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{`RANDOM}};
  _T_1013_im = _RAND_1651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{`RANDOM}};
  _T_1014_re = _RAND_1652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{`RANDOM}};
  _T_1014_im = _RAND_1653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{`RANDOM}};
  _T_1015_re = _RAND_1654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{`RANDOM}};
  _T_1015_im = _RAND_1655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{`RANDOM}};
  _T_1016_re = _RAND_1656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{`RANDOM}};
  _T_1016_im = _RAND_1657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{`RANDOM}};
  _T_1017_re = _RAND_1658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{`RANDOM}};
  _T_1017_im = _RAND_1659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{`RANDOM}};
  _T_1018_re = _RAND_1660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{`RANDOM}};
  _T_1018_im = _RAND_1661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{`RANDOM}};
  _T_1019_re = _RAND_1662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{`RANDOM}};
  _T_1019_im = _RAND_1663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{`RANDOM}};
  _T_1020_re = _RAND_1664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{`RANDOM}};
  _T_1020_im = _RAND_1665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{`RANDOM}};
  _T_1021_re = _RAND_1666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{`RANDOM}};
  _T_1021_im = _RAND_1667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{`RANDOM}};
  _T_1022_re = _RAND_1668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{`RANDOM}};
  _T_1022_im = _RAND_1669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{`RANDOM}};
  _T_1023_re = _RAND_1670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{`RANDOM}};
  _T_1023_im = _RAND_1671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{`RANDOM}};
  _T_1024_re = _RAND_1672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{`RANDOM}};
  _T_1024_im = _RAND_1673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{`RANDOM}};
  _T_1025_re = _RAND_1674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{`RANDOM}};
  _T_1025_im = _RAND_1675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{`RANDOM}};
  _T_1026_re = _RAND_1676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{`RANDOM}};
  _T_1026_im = _RAND_1677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{`RANDOM}};
  _T_1027_re = _RAND_1678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{`RANDOM}};
  _T_1027_im = _RAND_1679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{`RANDOM}};
  _T_1028_re = _RAND_1680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{`RANDOM}};
  _T_1028_im = _RAND_1681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{`RANDOM}};
  _T_1029_re = _RAND_1682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{`RANDOM}};
  _T_1029_im = _RAND_1683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{`RANDOM}};
  _T_1030_re = _RAND_1684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{`RANDOM}};
  _T_1030_im = _RAND_1685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{`RANDOM}};
  _T_1031_re = _RAND_1686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{`RANDOM}};
  _T_1031_im = _RAND_1687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{`RANDOM}};
  _T_1032_re = _RAND_1688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{`RANDOM}};
  _T_1032_im = _RAND_1689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{`RANDOM}};
  _T_1033_re = _RAND_1690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{`RANDOM}};
  _T_1033_im = _RAND_1691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{`RANDOM}};
  _T_1034_re = _RAND_1692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{`RANDOM}};
  _T_1034_im = _RAND_1693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{`RANDOM}};
  _T_1035_re = _RAND_1694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{`RANDOM}};
  _T_1035_im = _RAND_1695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{`RANDOM}};
  _T_1036_re = _RAND_1696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{`RANDOM}};
  _T_1036_im = _RAND_1697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{`RANDOM}};
  _T_1037_re = _RAND_1698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{`RANDOM}};
  _T_1037_im = _RAND_1699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{`RANDOM}};
  _T_1038_re = _RAND_1700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{`RANDOM}};
  _T_1038_im = _RAND_1701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{`RANDOM}};
  _T_1039_re = _RAND_1702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{`RANDOM}};
  _T_1039_im = _RAND_1703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{`RANDOM}};
  _T_1040_re = _RAND_1704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{`RANDOM}};
  _T_1040_im = _RAND_1705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{`RANDOM}};
  _T_1041_re = _RAND_1706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{`RANDOM}};
  _T_1041_im = _RAND_1707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{`RANDOM}};
  _T_1042_re = _RAND_1708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{`RANDOM}};
  _T_1042_im = _RAND_1709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{`RANDOM}};
  _T_1043_re = _RAND_1710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{`RANDOM}};
  _T_1043_im = _RAND_1711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{`RANDOM}};
  _T_1044_re = _RAND_1712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{`RANDOM}};
  _T_1044_im = _RAND_1713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{`RANDOM}};
  _T_1045_re = _RAND_1714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{`RANDOM}};
  _T_1045_im = _RAND_1715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{`RANDOM}};
  _T_1046_re = _RAND_1716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{`RANDOM}};
  _T_1046_im = _RAND_1717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{`RANDOM}};
  _T_1047_re = _RAND_1718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{`RANDOM}};
  _T_1047_im = _RAND_1719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{`RANDOM}};
  _T_1048_re = _RAND_1720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{`RANDOM}};
  _T_1048_im = _RAND_1721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{`RANDOM}};
  _T_1049_re = _RAND_1722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{`RANDOM}};
  _T_1049_im = _RAND_1723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{`RANDOM}};
  _T_1050_re = _RAND_1724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{`RANDOM}};
  _T_1050_im = _RAND_1725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{`RANDOM}};
  _T_1051_re = _RAND_1726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{`RANDOM}};
  _T_1051_im = _RAND_1727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{`RANDOM}};
  _T_1052_re = _RAND_1728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{`RANDOM}};
  _T_1052_im = _RAND_1729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{`RANDOM}};
  _T_1053_re = _RAND_1730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{`RANDOM}};
  _T_1053_im = _RAND_1731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{`RANDOM}};
  _T_1054_re = _RAND_1732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{`RANDOM}};
  _T_1054_im = _RAND_1733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{`RANDOM}};
  _T_1055_re = _RAND_1734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{`RANDOM}};
  _T_1055_im = _RAND_1735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{`RANDOM}};
  _T_1056_re = _RAND_1736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{`RANDOM}};
  _T_1056_im = _RAND_1737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{`RANDOM}};
  _T_1057_re = _RAND_1738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{`RANDOM}};
  _T_1057_im = _RAND_1739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{`RANDOM}};
  _T_1058_re = _RAND_1740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{`RANDOM}};
  _T_1058_im = _RAND_1741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{`RANDOM}};
  _T_1059_re = _RAND_1742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{`RANDOM}};
  _T_1059_im = _RAND_1743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{`RANDOM}};
  _T_1060_re = _RAND_1744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{`RANDOM}};
  _T_1060_im = _RAND_1745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{`RANDOM}};
  _T_1061_re = _RAND_1746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{`RANDOM}};
  _T_1061_im = _RAND_1747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{`RANDOM}};
  _T_1062_re = _RAND_1748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{`RANDOM}};
  _T_1062_im = _RAND_1749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{`RANDOM}};
  _T_1063_re = _RAND_1750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{`RANDOM}};
  _T_1063_im = _RAND_1751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{`RANDOM}};
  _T_1064_re = _RAND_1752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{`RANDOM}};
  _T_1064_im = _RAND_1753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{`RANDOM}};
  _T_1065_re = _RAND_1754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{`RANDOM}};
  _T_1065_im = _RAND_1755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{`RANDOM}};
  _T_1066_re = _RAND_1756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{`RANDOM}};
  _T_1066_im = _RAND_1757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{`RANDOM}};
  _T_1067_re = _RAND_1758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{`RANDOM}};
  _T_1067_im = _RAND_1759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{`RANDOM}};
  _T_1068_re = _RAND_1760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{`RANDOM}};
  _T_1068_im = _RAND_1761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{`RANDOM}};
  _T_1069_re = _RAND_1762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{`RANDOM}};
  _T_1069_im = _RAND_1763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{`RANDOM}};
  _T_1070_re = _RAND_1764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{`RANDOM}};
  _T_1070_im = _RAND_1765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{`RANDOM}};
  _T_1071_re = _RAND_1766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{`RANDOM}};
  _T_1071_im = _RAND_1767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{`RANDOM}};
  _T_1072_re = _RAND_1768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{`RANDOM}};
  _T_1072_im = _RAND_1769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{`RANDOM}};
  _T_1073_re = _RAND_1770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{`RANDOM}};
  _T_1073_im = _RAND_1771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{`RANDOM}};
  _T_1074_re = _RAND_1772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{`RANDOM}};
  _T_1074_im = _RAND_1773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{`RANDOM}};
  _T_1075_re = _RAND_1774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{`RANDOM}};
  _T_1075_im = _RAND_1775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{`RANDOM}};
  _T_1076_re = _RAND_1776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{`RANDOM}};
  _T_1076_im = _RAND_1777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{`RANDOM}};
  _T_1077_re = _RAND_1778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{`RANDOM}};
  _T_1077_im = _RAND_1779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{`RANDOM}};
  _T_1078_re = _RAND_1780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{`RANDOM}};
  _T_1078_im = _RAND_1781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{`RANDOM}};
  _T_1079_re = _RAND_1782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{`RANDOM}};
  _T_1079_im = _RAND_1783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{`RANDOM}};
  _T_1080_re = _RAND_1784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{`RANDOM}};
  _T_1080_im = _RAND_1785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{`RANDOM}};
  _T_1081_re = _RAND_1786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{`RANDOM}};
  _T_1081_im = _RAND_1787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{`RANDOM}};
  _T_1082_re = _RAND_1788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{`RANDOM}};
  _T_1082_im = _RAND_1789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{`RANDOM}};
  _T_1083_re = _RAND_1790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{`RANDOM}};
  _T_1083_im = _RAND_1791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{`RANDOM}};
  _T_1084_re = _RAND_1792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{`RANDOM}};
  _T_1084_im = _RAND_1793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{`RANDOM}};
  _T_1085_re = _RAND_1794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{`RANDOM}};
  _T_1085_im = _RAND_1795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{`RANDOM}};
  _T_1086_re = _RAND_1796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{`RANDOM}};
  _T_1086_im = _RAND_1797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{`RANDOM}};
  _T_1087_re = _RAND_1798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{`RANDOM}};
  _T_1087_im = _RAND_1799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{`RANDOM}};
  _T_1088_re = _RAND_1800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{`RANDOM}};
  _T_1088_im = _RAND_1801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{`RANDOM}};
  _T_1089_re = _RAND_1802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{`RANDOM}};
  _T_1089_im = _RAND_1803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{`RANDOM}};
  _T_1090_re = _RAND_1804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{`RANDOM}};
  _T_1090_im = _RAND_1805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{`RANDOM}};
  _T_1091_re = _RAND_1806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{`RANDOM}};
  _T_1091_im = _RAND_1807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{`RANDOM}};
  _T_1092_re = _RAND_1808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{`RANDOM}};
  _T_1092_im = _RAND_1809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{`RANDOM}};
  _T_1093_re = _RAND_1810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{`RANDOM}};
  _T_1093_im = _RAND_1811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{`RANDOM}};
  _T_1094_re = _RAND_1812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{`RANDOM}};
  _T_1094_im = _RAND_1813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{`RANDOM}};
  _T_1095_re = _RAND_1814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{`RANDOM}};
  _T_1095_im = _RAND_1815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{`RANDOM}};
  _T_1096_re = _RAND_1816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{`RANDOM}};
  _T_1096_im = _RAND_1817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{`RANDOM}};
  _T_1097_re = _RAND_1818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{`RANDOM}};
  _T_1097_im = _RAND_1819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{`RANDOM}};
  _T_1098_re = _RAND_1820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{`RANDOM}};
  _T_1098_im = _RAND_1821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{`RANDOM}};
  _T_1099_re = _RAND_1822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{`RANDOM}};
  _T_1099_im = _RAND_1823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{`RANDOM}};
  _T_1100_re = _RAND_1824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{`RANDOM}};
  _T_1100_im = _RAND_1825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{`RANDOM}};
  _T_1101_re = _RAND_1826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{`RANDOM}};
  _T_1101_im = _RAND_1827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{`RANDOM}};
  _T_1102_re = _RAND_1828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{`RANDOM}};
  _T_1102_im = _RAND_1829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{`RANDOM}};
  _T_1103_re = _RAND_1830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{`RANDOM}};
  _T_1103_im = _RAND_1831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{`RANDOM}};
  _T_1104_re = _RAND_1832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{`RANDOM}};
  _T_1104_im = _RAND_1833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{`RANDOM}};
  _T_1105_re = _RAND_1834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{`RANDOM}};
  _T_1105_im = _RAND_1835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{`RANDOM}};
  _T_1106_re = _RAND_1836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{`RANDOM}};
  _T_1106_im = _RAND_1837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{`RANDOM}};
  _T_1107_re = _RAND_1838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{`RANDOM}};
  _T_1107_im = _RAND_1839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{`RANDOM}};
  _T_1108_re = _RAND_1840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{`RANDOM}};
  _T_1108_im = _RAND_1841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{`RANDOM}};
  _T_1109_re = _RAND_1842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{`RANDOM}};
  _T_1109_im = _RAND_1843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{`RANDOM}};
  _T_1110_re = _RAND_1844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{`RANDOM}};
  _T_1110_im = _RAND_1845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{`RANDOM}};
  _T_1111_re = _RAND_1846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{`RANDOM}};
  _T_1111_im = _RAND_1847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{`RANDOM}};
  _T_1112_re = _RAND_1848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{`RANDOM}};
  _T_1112_im = _RAND_1849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{`RANDOM}};
  _T_1113_re = _RAND_1850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{`RANDOM}};
  _T_1113_im = _RAND_1851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{`RANDOM}};
  _T_1114_re = _RAND_1852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{`RANDOM}};
  _T_1114_im = _RAND_1853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{`RANDOM}};
  _T_1115_re = _RAND_1854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{`RANDOM}};
  _T_1115_im = _RAND_1855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{`RANDOM}};
  _T_1116_re = _RAND_1856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{`RANDOM}};
  _T_1116_im = _RAND_1857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{`RANDOM}};
  _T_1117_re = _RAND_1858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{`RANDOM}};
  _T_1117_im = _RAND_1859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{`RANDOM}};
  _T_1118_re = _RAND_1860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{`RANDOM}};
  _T_1118_im = _RAND_1861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{`RANDOM}};
  _T_1119_re = _RAND_1862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{`RANDOM}};
  _T_1119_im = _RAND_1863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{`RANDOM}};
  _T_1120_re = _RAND_1864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{`RANDOM}};
  _T_1120_im = _RAND_1865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{`RANDOM}};
  _T_1121_re = _RAND_1866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{`RANDOM}};
  _T_1121_im = _RAND_1867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{`RANDOM}};
  _T_1122_re = _RAND_1868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{`RANDOM}};
  _T_1122_im = _RAND_1869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{`RANDOM}};
  _T_1123_re = _RAND_1870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{`RANDOM}};
  _T_1123_im = _RAND_1871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{`RANDOM}};
  _T_1124_re = _RAND_1872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{`RANDOM}};
  _T_1124_im = _RAND_1873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{`RANDOM}};
  _T_1125_re = _RAND_1874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{`RANDOM}};
  _T_1125_im = _RAND_1875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{`RANDOM}};
  _T_1126_re = _RAND_1876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{`RANDOM}};
  _T_1126_im = _RAND_1877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{`RANDOM}};
  _T_1127_re = _RAND_1878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{`RANDOM}};
  _T_1127_im = _RAND_1879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{`RANDOM}};
  _T_1128_re = _RAND_1880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{`RANDOM}};
  _T_1128_im = _RAND_1881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{`RANDOM}};
  _T_1129_re = _RAND_1882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{`RANDOM}};
  _T_1129_im = _RAND_1883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{`RANDOM}};
  _T_1130_re = _RAND_1884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{`RANDOM}};
  _T_1130_im = _RAND_1885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{`RANDOM}};
  _T_1131_re = _RAND_1886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{`RANDOM}};
  _T_1131_im = _RAND_1887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{`RANDOM}};
  _T_1132_re = _RAND_1888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{`RANDOM}};
  _T_1132_im = _RAND_1889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{`RANDOM}};
  _T_1133_re = _RAND_1890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{`RANDOM}};
  _T_1133_im = _RAND_1891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{`RANDOM}};
  _T_1134_re = _RAND_1892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{`RANDOM}};
  _T_1134_im = _RAND_1893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{`RANDOM}};
  _T_1135_re = _RAND_1894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{`RANDOM}};
  _T_1135_im = _RAND_1895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{`RANDOM}};
  _T_1136_re = _RAND_1896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{`RANDOM}};
  _T_1136_im = _RAND_1897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{`RANDOM}};
  _T_1137_re = _RAND_1898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{`RANDOM}};
  _T_1137_im = _RAND_1899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{`RANDOM}};
  _T_1138_re = _RAND_1900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{`RANDOM}};
  _T_1138_im = _RAND_1901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{`RANDOM}};
  _T_1139_re = _RAND_1902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{`RANDOM}};
  _T_1139_im = _RAND_1903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{`RANDOM}};
  _T_1140_re = _RAND_1904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{`RANDOM}};
  _T_1140_im = _RAND_1905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{`RANDOM}};
  _T_1141_re = _RAND_1906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{`RANDOM}};
  _T_1141_im = _RAND_1907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{`RANDOM}};
  _T_1142_re = _RAND_1908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{`RANDOM}};
  _T_1142_im = _RAND_1909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{`RANDOM}};
  _T_1143_re = _RAND_1910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{`RANDOM}};
  _T_1143_im = _RAND_1911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{`RANDOM}};
  _T_1144_re = _RAND_1912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{`RANDOM}};
  _T_1144_im = _RAND_1913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{`RANDOM}};
  _T_1145_re = _RAND_1914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{`RANDOM}};
  _T_1145_im = _RAND_1915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{`RANDOM}};
  _T_1146_re = _RAND_1916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{`RANDOM}};
  _T_1146_im = _RAND_1917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{`RANDOM}};
  _T_1147_re = _RAND_1918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{`RANDOM}};
  _T_1147_im = _RAND_1919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{`RANDOM}};
  _T_1148_re = _RAND_1920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{`RANDOM}};
  _T_1148_im = _RAND_1921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{`RANDOM}};
  _T_1149_re = _RAND_1922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{`RANDOM}};
  _T_1149_im = _RAND_1923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{`RANDOM}};
  _T_1150_re = _RAND_1924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{`RANDOM}};
  _T_1150_im = _RAND_1925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{`RANDOM}};
  _T_1151_re = _RAND_1926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{`RANDOM}};
  _T_1151_im = _RAND_1927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{`RANDOM}};
  _T_1152_re = _RAND_1928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{`RANDOM}};
  _T_1152_im = _RAND_1929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{`RANDOM}};
  _T_1153_re = _RAND_1930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{`RANDOM}};
  _T_1153_im = _RAND_1931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{`RANDOM}};
  _T_1154_re = _RAND_1932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{`RANDOM}};
  _T_1154_im = _RAND_1933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{`RANDOM}};
  _T_1155_re = _RAND_1934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{`RANDOM}};
  _T_1155_im = _RAND_1935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{`RANDOM}};
  _T_1156_re = _RAND_1936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{`RANDOM}};
  _T_1156_im = _RAND_1937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{`RANDOM}};
  _T_1157_re = _RAND_1938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{`RANDOM}};
  _T_1157_im = _RAND_1939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{`RANDOM}};
  _T_1158_re = _RAND_1940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{`RANDOM}};
  _T_1158_im = _RAND_1941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{`RANDOM}};
  _T_1159_re = _RAND_1942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{`RANDOM}};
  _T_1159_im = _RAND_1943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{`RANDOM}};
  _T_1160_re = _RAND_1944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{`RANDOM}};
  _T_1160_im = _RAND_1945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{`RANDOM}};
  _T_1161_re = _RAND_1946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{`RANDOM}};
  _T_1161_im = _RAND_1947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{`RANDOM}};
  _T_1162_re = _RAND_1948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{`RANDOM}};
  _T_1162_im = _RAND_1949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{`RANDOM}};
  _T_1163_re = _RAND_1950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{`RANDOM}};
  _T_1163_im = _RAND_1951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{`RANDOM}};
  _T_1164_re = _RAND_1952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{`RANDOM}};
  _T_1164_im = _RAND_1953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{`RANDOM}};
  _T_1165_re = _RAND_1954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{`RANDOM}};
  _T_1165_im = _RAND_1955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{`RANDOM}};
  _T_1166_re = _RAND_1956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{`RANDOM}};
  _T_1166_im = _RAND_1957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{`RANDOM}};
  _T_1167_re = _RAND_1958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{`RANDOM}};
  _T_1167_im = _RAND_1959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{`RANDOM}};
  _T_1168_re = _RAND_1960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{`RANDOM}};
  _T_1168_im = _RAND_1961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{`RANDOM}};
  _T_1169_re = _RAND_1962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{`RANDOM}};
  _T_1169_im = _RAND_1963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{`RANDOM}};
  _T_1170_re = _RAND_1964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{`RANDOM}};
  _T_1170_im = _RAND_1965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{`RANDOM}};
  _T_1171_re = _RAND_1966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{`RANDOM}};
  _T_1171_im = _RAND_1967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{`RANDOM}};
  _T_1172_re = _RAND_1968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{`RANDOM}};
  _T_1172_im = _RAND_1969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{`RANDOM}};
  _T_1173_re = _RAND_1970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{`RANDOM}};
  _T_1173_im = _RAND_1971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{`RANDOM}};
  _T_1174_re = _RAND_1972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{`RANDOM}};
  _T_1174_im = _RAND_1973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{`RANDOM}};
  _T_1175_re = _RAND_1974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{`RANDOM}};
  _T_1175_im = _RAND_1975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{`RANDOM}};
  _T_1176_re = _RAND_1976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{`RANDOM}};
  _T_1176_im = _RAND_1977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{`RANDOM}};
  _T_1177_re = _RAND_1978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{`RANDOM}};
  _T_1177_im = _RAND_1979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{`RANDOM}};
  _T_1178_re = _RAND_1980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{`RANDOM}};
  _T_1178_im = _RAND_1981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{`RANDOM}};
  _T_1179_re = _RAND_1982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{`RANDOM}};
  _T_1179_im = _RAND_1983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{`RANDOM}};
  _T_1180_re = _RAND_1984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{`RANDOM}};
  _T_1180_im = _RAND_1985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{`RANDOM}};
  _T_1181_re = _RAND_1986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{`RANDOM}};
  _T_1181_im = _RAND_1987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{`RANDOM}};
  _T_1182_re = _RAND_1988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{`RANDOM}};
  _T_1182_im = _RAND_1989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{`RANDOM}};
  _T_1183_re = _RAND_1990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{`RANDOM}};
  _T_1183_im = _RAND_1991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{`RANDOM}};
  _T_1184_re = _RAND_1992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{`RANDOM}};
  _T_1184_im = _RAND_1993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{`RANDOM}};
  _T_1185_re = _RAND_1994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{`RANDOM}};
  _T_1185_im = _RAND_1995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{`RANDOM}};
  _T_1186_re = _RAND_1996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{`RANDOM}};
  _T_1186_im = _RAND_1997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{`RANDOM}};
  _T_1187_re = _RAND_1998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{`RANDOM}};
  _T_1187_im = _RAND_1999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{`RANDOM}};
  _T_1188_re = _RAND_2000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{`RANDOM}};
  _T_1188_im = _RAND_2001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{`RANDOM}};
  _T_1189_re = _RAND_2002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{`RANDOM}};
  _T_1189_im = _RAND_2003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{`RANDOM}};
  _T_1190_re = _RAND_2004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{`RANDOM}};
  _T_1190_im = _RAND_2005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{`RANDOM}};
  _T_1191_re = _RAND_2006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{`RANDOM}};
  _T_1191_im = _RAND_2007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{`RANDOM}};
  _T_1192_re = _RAND_2008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{`RANDOM}};
  _T_1192_im = _RAND_2009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{`RANDOM}};
  _T_1193_re = _RAND_2010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{`RANDOM}};
  _T_1193_im = _RAND_2011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{`RANDOM}};
  _T_1194_re = _RAND_2012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{`RANDOM}};
  _T_1194_im = _RAND_2013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{`RANDOM}};
  _T_1195_re = _RAND_2014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{`RANDOM}};
  _T_1195_im = _RAND_2015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{`RANDOM}};
  _T_1196_re = _RAND_2016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{`RANDOM}};
  _T_1196_im = _RAND_2017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{`RANDOM}};
  _T_1197_re = _RAND_2018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{`RANDOM}};
  _T_1197_im = _RAND_2019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{`RANDOM}};
  _T_1198_re = _RAND_2020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{`RANDOM}};
  _T_1198_im = _RAND_2021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{`RANDOM}};
  _T_1199_re = _RAND_2022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{`RANDOM}};
  _T_1199_im = _RAND_2023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{`RANDOM}};
  _T_1200_re = _RAND_2024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{`RANDOM}};
  _T_1200_im = _RAND_2025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{`RANDOM}};
  _T_1201_re = _RAND_2026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{`RANDOM}};
  _T_1201_im = _RAND_2027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{`RANDOM}};
  _T_1202_re = _RAND_2028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{`RANDOM}};
  _T_1202_im = _RAND_2029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{`RANDOM}};
  _T_1203_re = _RAND_2030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{`RANDOM}};
  _T_1203_im = _RAND_2031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{`RANDOM}};
  _T_1204_re = _RAND_2032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{`RANDOM}};
  _T_1204_im = _RAND_2033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{`RANDOM}};
  _T_1205_re = _RAND_2034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{`RANDOM}};
  _T_1205_im = _RAND_2035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{`RANDOM}};
  _T_1206_re = _RAND_2036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{`RANDOM}};
  _T_1206_im = _RAND_2037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{`RANDOM}};
  _T_1207_re = _RAND_2038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{`RANDOM}};
  _T_1207_im = _RAND_2039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{`RANDOM}};
  _T_1208_re = _RAND_2040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{`RANDOM}};
  _T_1208_im = _RAND_2041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{`RANDOM}};
  _T_1209_re = _RAND_2042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{`RANDOM}};
  _T_1209_im = _RAND_2043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{`RANDOM}};
  _T_1210_re = _RAND_2044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{`RANDOM}};
  _T_1210_im = _RAND_2045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{`RANDOM}};
  _T_1211_re = _RAND_2046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{`RANDOM}};
  _T_1211_im = _RAND_2047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2048 = {1{`RANDOM}};
  _T_1212_re = _RAND_2048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2049 = {1{`RANDOM}};
  _T_1212_im = _RAND_2049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2050 = {1{`RANDOM}};
  _T_1213_re = _RAND_2050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2051 = {1{`RANDOM}};
  _T_1213_im = _RAND_2051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2052 = {1{`RANDOM}};
  _T_1214_re = _RAND_2052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2053 = {1{`RANDOM}};
  _T_1214_im = _RAND_2053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2054 = {1{`RANDOM}};
  _T_1215_re = _RAND_2054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2055 = {1{`RANDOM}};
  _T_1215_im = _RAND_2055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2056 = {1{`RANDOM}};
  _T_1216_re = _RAND_2056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2057 = {1{`RANDOM}};
  _T_1216_im = _RAND_2057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2058 = {1{`RANDOM}};
  _T_1217_re = _RAND_2058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2059 = {1{`RANDOM}};
  _T_1217_im = _RAND_2059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2060 = {1{`RANDOM}};
  _T_1218_re = _RAND_2060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2061 = {1{`RANDOM}};
  _T_1218_im = _RAND_2061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2062 = {1{`RANDOM}};
  _T_1219_re = _RAND_2062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2063 = {1{`RANDOM}};
  _T_1219_im = _RAND_2063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2064 = {1{`RANDOM}};
  _T_1220_re = _RAND_2064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2065 = {1{`RANDOM}};
  _T_1220_im = _RAND_2065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2066 = {1{`RANDOM}};
  _T_1221_re = _RAND_2066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2067 = {1{`RANDOM}};
  _T_1221_im = _RAND_2067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2068 = {1{`RANDOM}};
  _T_1222_re = _RAND_2068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2069 = {1{`RANDOM}};
  _T_1222_im = _RAND_2069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2070 = {1{`RANDOM}};
  _T_1223_re = _RAND_2070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2071 = {1{`RANDOM}};
  _T_1223_im = _RAND_2071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2072 = {1{`RANDOM}};
  _T_1224_re = _RAND_2072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2073 = {1{`RANDOM}};
  _T_1224_im = _RAND_2073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2074 = {1{`RANDOM}};
  _T_1225_re = _RAND_2074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2075 = {1{`RANDOM}};
  _T_1225_im = _RAND_2075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2076 = {1{`RANDOM}};
  _T_1226_re = _RAND_2076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2077 = {1{`RANDOM}};
  _T_1226_im = _RAND_2077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2078 = {1{`RANDOM}};
  _T_1227_re = _RAND_2078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2079 = {1{`RANDOM}};
  _T_1227_im = _RAND_2079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2080 = {1{`RANDOM}};
  _T_1228_re = _RAND_2080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2081 = {1{`RANDOM}};
  _T_1228_im = _RAND_2081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2082 = {1{`RANDOM}};
  _T_1229_re = _RAND_2082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2083 = {1{`RANDOM}};
  _T_1229_im = _RAND_2083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2084 = {1{`RANDOM}};
  _T_1230_re = _RAND_2084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2085 = {1{`RANDOM}};
  _T_1230_im = _RAND_2085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2086 = {1{`RANDOM}};
  _T_1231_re = _RAND_2086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2087 = {1{`RANDOM}};
  _T_1231_im = _RAND_2087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2088 = {1{`RANDOM}};
  _T_1232_re = _RAND_2088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2089 = {1{`RANDOM}};
  _T_1232_im = _RAND_2089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2090 = {1{`RANDOM}};
  _T_1233_re = _RAND_2090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2091 = {1{`RANDOM}};
  _T_1233_im = _RAND_2091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2092 = {1{`RANDOM}};
  _T_1234_re = _RAND_2092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2093 = {1{`RANDOM}};
  _T_1234_im = _RAND_2093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2094 = {1{`RANDOM}};
  _T_1235_re = _RAND_2094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2095 = {1{`RANDOM}};
  _T_1235_im = _RAND_2095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2096 = {1{`RANDOM}};
  _T_1236_re = _RAND_2096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2097 = {1{`RANDOM}};
  _T_1236_im = _RAND_2097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2098 = {1{`RANDOM}};
  _T_1237_re = _RAND_2098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2099 = {1{`RANDOM}};
  _T_1237_im = _RAND_2099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2100 = {1{`RANDOM}};
  _T_1238_re = _RAND_2100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2101 = {1{`RANDOM}};
  _T_1238_im = _RAND_2101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2102 = {1{`RANDOM}};
  _T_1239_re = _RAND_2102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2103 = {1{`RANDOM}};
  _T_1239_im = _RAND_2103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2104 = {1{`RANDOM}};
  _T_1240_re = _RAND_2104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2105 = {1{`RANDOM}};
  _T_1240_im = _RAND_2105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2106 = {1{`RANDOM}};
  _T_1241_re = _RAND_2106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2107 = {1{`RANDOM}};
  _T_1241_im = _RAND_2107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2108 = {1{`RANDOM}};
  _T_1242_re = _RAND_2108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2109 = {1{`RANDOM}};
  _T_1242_im = _RAND_2109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2110 = {1{`RANDOM}};
  _T_1243_re = _RAND_2110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2111 = {1{`RANDOM}};
  _T_1243_im = _RAND_2111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2112 = {1{`RANDOM}};
  _T_1244_re = _RAND_2112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2113 = {1{`RANDOM}};
  _T_1244_im = _RAND_2113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2114 = {1{`RANDOM}};
  _T_1245_re = _RAND_2114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2115 = {1{`RANDOM}};
  _T_1245_im = _RAND_2115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2116 = {1{`RANDOM}};
  _T_1246_re = _RAND_2116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2117 = {1{`RANDOM}};
  _T_1246_im = _RAND_2117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2118 = {1{`RANDOM}};
  _T_1247_re = _RAND_2118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2119 = {1{`RANDOM}};
  _T_1247_im = _RAND_2119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2120 = {1{`RANDOM}};
  _T_1248_re = _RAND_2120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2121 = {1{`RANDOM}};
  _T_1248_im = _RAND_2121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2122 = {1{`RANDOM}};
  _T_1249_re = _RAND_2122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2123 = {1{`RANDOM}};
  _T_1249_im = _RAND_2123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2124 = {1{`RANDOM}};
  _T_1250_re = _RAND_2124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2125 = {1{`RANDOM}};
  _T_1250_im = _RAND_2125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2126 = {1{`RANDOM}};
  _T_1251_re = _RAND_2126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2127 = {1{`RANDOM}};
  _T_1251_im = _RAND_2127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2128 = {1{`RANDOM}};
  _T_1252_re = _RAND_2128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2129 = {1{`RANDOM}};
  _T_1252_im = _RAND_2129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2130 = {1{`RANDOM}};
  _T_1253_re = _RAND_2130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2131 = {1{`RANDOM}};
  _T_1253_im = _RAND_2131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2132 = {1{`RANDOM}};
  _T_1254_re = _RAND_2132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2133 = {1{`RANDOM}};
  _T_1254_im = _RAND_2133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2134 = {1{`RANDOM}};
  _T_1255_re = _RAND_2134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2135 = {1{`RANDOM}};
  _T_1255_im = _RAND_2135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2136 = {1{`RANDOM}};
  _T_1256_re = _RAND_2136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2137 = {1{`RANDOM}};
  _T_1256_im = _RAND_2137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2138 = {1{`RANDOM}};
  _T_1257_re = _RAND_2138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2139 = {1{`RANDOM}};
  _T_1257_im = _RAND_2139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2140 = {1{`RANDOM}};
  _T_1258_re = _RAND_2140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2141 = {1{`RANDOM}};
  _T_1258_im = _RAND_2141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2142 = {1{`RANDOM}};
  _T_1259_re = _RAND_2142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2143 = {1{`RANDOM}};
  _T_1259_im = _RAND_2143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2144 = {1{`RANDOM}};
  _T_1260_re = _RAND_2144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2145 = {1{`RANDOM}};
  _T_1260_im = _RAND_2145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2146 = {1{`RANDOM}};
  _T_1261_re = _RAND_2146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2147 = {1{`RANDOM}};
  _T_1261_im = _RAND_2147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2148 = {1{`RANDOM}};
  _T_1262_re = _RAND_2148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2149 = {1{`RANDOM}};
  _T_1262_im = _RAND_2149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2150 = {1{`RANDOM}};
  _T_1263_re = _RAND_2150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2151 = {1{`RANDOM}};
  _T_1263_im = _RAND_2151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2152 = {1{`RANDOM}};
  _T_1264_re = _RAND_2152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2153 = {1{`RANDOM}};
  _T_1264_im = _RAND_2153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2154 = {1{`RANDOM}};
  _T_1265_re = _RAND_2154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2155 = {1{`RANDOM}};
  _T_1265_im = _RAND_2155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2156 = {1{`RANDOM}};
  _T_1266_re = _RAND_2156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2157 = {1{`RANDOM}};
  _T_1266_im = _RAND_2157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2158 = {1{`RANDOM}};
  _T_1267_re = _RAND_2158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2159 = {1{`RANDOM}};
  _T_1267_im = _RAND_2159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2160 = {1{`RANDOM}};
  _T_1268_re = _RAND_2160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2161 = {1{`RANDOM}};
  _T_1268_im = _RAND_2161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2162 = {1{`RANDOM}};
  _T_1269_re = _RAND_2162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2163 = {1{`RANDOM}};
  _T_1269_im = _RAND_2163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2164 = {1{`RANDOM}};
  _T_1270_re = _RAND_2164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2165 = {1{`RANDOM}};
  _T_1270_im = _RAND_2165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2166 = {1{`RANDOM}};
  _T_1271_re = _RAND_2166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2167 = {1{`RANDOM}};
  _T_1271_im = _RAND_2167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2168 = {1{`RANDOM}};
  _T_1272_re = _RAND_2168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2169 = {1{`RANDOM}};
  _T_1272_im = _RAND_2169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2170 = {1{`RANDOM}};
  _T_1273_re = _RAND_2170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2171 = {1{`RANDOM}};
  _T_1273_im = _RAND_2171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2172 = {1{`RANDOM}};
  _T_1274_re = _RAND_2172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2173 = {1{`RANDOM}};
  _T_1274_im = _RAND_2173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2174 = {1{`RANDOM}};
  _T_1275_re = _RAND_2174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2175 = {1{`RANDOM}};
  _T_1275_im = _RAND_2175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2176 = {1{`RANDOM}};
  _T_1276_re = _RAND_2176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2177 = {1{`RANDOM}};
  _T_1276_im = _RAND_2177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2178 = {1{`RANDOM}};
  _T_1277_re = _RAND_2178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2179 = {1{`RANDOM}};
  _T_1277_im = _RAND_2179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2180 = {1{`RANDOM}};
  _T_1278_re = _RAND_2180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2181 = {1{`RANDOM}};
  _T_1278_im = _RAND_2181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2182 = {1{`RANDOM}};
  _T_1279_re = _RAND_2182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2183 = {1{`RANDOM}};
  _T_1279_im = _RAND_2183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2184 = {1{`RANDOM}};
  _T_1280_re = _RAND_2184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2185 = {1{`RANDOM}};
  _T_1280_im = _RAND_2185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2186 = {1{`RANDOM}};
  _T_1281_re = _RAND_2186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2187 = {1{`RANDOM}};
  _T_1281_im = _RAND_2187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2188 = {1{`RANDOM}};
  _T_1282_re = _RAND_2188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2189 = {1{`RANDOM}};
  _T_1282_im = _RAND_2189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2190 = {1{`RANDOM}};
  _T_1283_re = _RAND_2190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2191 = {1{`RANDOM}};
  _T_1283_im = _RAND_2191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2192 = {1{`RANDOM}};
  _T_1284_re = _RAND_2192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2193 = {1{`RANDOM}};
  _T_1284_im = _RAND_2193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2194 = {1{`RANDOM}};
  _T_1285_re = _RAND_2194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2195 = {1{`RANDOM}};
  _T_1285_im = _RAND_2195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2196 = {1{`RANDOM}};
  _T_1286_re = _RAND_2196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2197 = {1{`RANDOM}};
  _T_1286_im = _RAND_2197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2198 = {1{`RANDOM}};
  _T_1287_re = _RAND_2198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2199 = {1{`RANDOM}};
  _T_1287_im = _RAND_2199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2200 = {1{`RANDOM}};
  _T_1288_re = _RAND_2200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2201 = {1{`RANDOM}};
  _T_1288_im = _RAND_2201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2202 = {1{`RANDOM}};
  _T_1289_re = _RAND_2202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2203 = {1{`RANDOM}};
  _T_1289_im = _RAND_2203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2204 = {1{`RANDOM}};
  _T_1290_re = _RAND_2204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2205 = {1{`RANDOM}};
  _T_1290_im = _RAND_2205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2206 = {1{`RANDOM}};
  _T_1291_re = _RAND_2206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2207 = {1{`RANDOM}};
  _T_1291_im = _RAND_2207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2208 = {1{`RANDOM}};
  _T_1292_re = _RAND_2208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2209 = {1{`RANDOM}};
  _T_1292_im = _RAND_2209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2210 = {1{`RANDOM}};
  _T_1293_re = _RAND_2210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2211 = {1{`RANDOM}};
  _T_1293_im = _RAND_2211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2212 = {1{`RANDOM}};
  _T_1294_re = _RAND_2212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2213 = {1{`RANDOM}};
  _T_1294_im = _RAND_2213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2214 = {1{`RANDOM}};
  _T_1295_re = _RAND_2214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2215 = {1{`RANDOM}};
  _T_1295_im = _RAND_2215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2216 = {1{`RANDOM}};
  _T_1296_re = _RAND_2216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2217 = {1{`RANDOM}};
  _T_1296_im = _RAND_2217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2218 = {1{`RANDOM}};
  _T_1297_re = _RAND_2218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2219 = {1{`RANDOM}};
  _T_1297_im = _RAND_2219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2220 = {1{`RANDOM}};
  _T_1298_re = _RAND_2220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2221 = {1{`RANDOM}};
  _T_1298_im = _RAND_2221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2222 = {1{`RANDOM}};
  _T_1299_re = _RAND_2222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2223 = {1{`RANDOM}};
  _T_1299_im = _RAND_2223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2224 = {1{`RANDOM}};
  _T_1300_re = _RAND_2224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2225 = {1{`RANDOM}};
  _T_1300_im = _RAND_2225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2226 = {1{`RANDOM}};
  _T_1301_re = _RAND_2226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2227 = {1{`RANDOM}};
  _T_1301_im = _RAND_2227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2228 = {1{`RANDOM}};
  _T_1302_re = _RAND_2228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2229 = {1{`RANDOM}};
  _T_1302_im = _RAND_2229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2230 = {1{`RANDOM}};
  _T_1303_re = _RAND_2230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2231 = {1{`RANDOM}};
  _T_1303_im = _RAND_2231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2232 = {1{`RANDOM}};
  _T_1304_re = _RAND_2232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2233 = {1{`RANDOM}};
  _T_1304_im = _RAND_2233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2234 = {1{`RANDOM}};
  _T_1305_re = _RAND_2234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2235 = {1{`RANDOM}};
  _T_1305_im = _RAND_2235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2236 = {1{`RANDOM}};
  _T_1306_re = _RAND_2236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2237 = {1{`RANDOM}};
  _T_1306_im = _RAND_2237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2238 = {1{`RANDOM}};
  _T_1307_re = _RAND_2238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2239 = {1{`RANDOM}};
  _T_1307_im = _RAND_2239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2240 = {1{`RANDOM}};
  _T_1308_re = _RAND_2240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2241 = {1{`RANDOM}};
  _T_1308_im = _RAND_2241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2242 = {1{`RANDOM}};
  _T_1309_re = _RAND_2242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2243 = {1{`RANDOM}};
  _T_1309_im = _RAND_2243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2244 = {1{`RANDOM}};
  _T_1310_re = _RAND_2244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2245 = {1{`RANDOM}};
  _T_1310_im = _RAND_2245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2246 = {1{`RANDOM}};
  _T_1311_re = _RAND_2246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2247 = {1{`RANDOM}};
  _T_1311_im = _RAND_2247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2248 = {1{`RANDOM}};
  _T_1312_re = _RAND_2248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2249 = {1{`RANDOM}};
  _T_1312_im = _RAND_2249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2250 = {1{`RANDOM}};
  _T_1313_re = _RAND_2250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2251 = {1{`RANDOM}};
  _T_1313_im = _RAND_2251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2252 = {1{`RANDOM}};
  _T_1314_re = _RAND_2252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2253 = {1{`RANDOM}};
  _T_1314_im = _RAND_2253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2254 = {1{`RANDOM}};
  _T_1315_re = _RAND_2254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2255 = {1{`RANDOM}};
  _T_1315_im = _RAND_2255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2256 = {1{`RANDOM}};
  _T_1316_re = _RAND_2256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2257 = {1{`RANDOM}};
  _T_1316_im = _RAND_2257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2258 = {1{`RANDOM}};
  _T_1317_re = _RAND_2258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2259 = {1{`RANDOM}};
  _T_1317_im = _RAND_2259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2260 = {1{`RANDOM}};
  _T_1318_re = _RAND_2260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2261 = {1{`RANDOM}};
  _T_1318_im = _RAND_2261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2262 = {1{`RANDOM}};
  _T_1319_re = _RAND_2262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2263 = {1{`RANDOM}};
  _T_1319_im = _RAND_2263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2264 = {1{`RANDOM}};
  _T_1320_re = _RAND_2264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2265 = {1{`RANDOM}};
  _T_1320_im = _RAND_2265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2266 = {1{`RANDOM}};
  _T_1321_re = _RAND_2266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2267 = {1{`RANDOM}};
  _T_1321_im = _RAND_2267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2268 = {1{`RANDOM}};
  _T_1322_re = _RAND_2268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2269 = {1{`RANDOM}};
  _T_1322_im = _RAND_2269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2270 = {1{`RANDOM}};
  _T_1323_re = _RAND_2270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2271 = {1{`RANDOM}};
  _T_1323_im = _RAND_2271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2272 = {1{`RANDOM}};
  _T_1324_re = _RAND_2272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2273 = {1{`RANDOM}};
  _T_1324_im = _RAND_2273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2274 = {1{`RANDOM}};
  _T_1325_re = _RAND_2274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2275 = {1{`RANDOM}};
  _T_1325_im = _RAND_2275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2276 = {1{`RANDOM}};
  _T_1326_re = _RAND_2276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2277 = {1{`RANDOM}};
  _T_1326_im = _RAND_2277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2278 = {1{`RANDOM}};
  _T_1327_re = _RAND_2278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2279 = {1{`RANDOM}};
  _T_1327_im = _RAND_2279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2280 = {1{`RANDOM}};
  _T_1328_re = _RAND_2280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2281 = {1{`RANDOM}};
  _T_1328_im = _RAND_2281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2282 = {1{`RANDOM}};
  _T_1329_re = _RAND_2282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2283 = {1{`RANDOM}};
  _T_1329_im = _RAND_2283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2284 = {1{`RANDOM}};
  _T_1330_re = _RAND_2284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2285 = {1{`RANDOM}};
  _T_1330_im = _RAND_2285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2286 = {1{`RANDOM}};
  _T_1331_re = _RAND_2286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2287 = {1{`RANDOM}};
  _T_1331_im = _RAND_2287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2288 = {1{`RANDOM}};
  _T_1332_re = _RAND_2288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2289 = {1{`RANDOM}};
  _T_1332_im = _RAND_2289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2290 = {1{`RANDOM}};
  _T_1333_re = _RAND_2290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2291 = {1{`RANDOM}};
  _T_1333_im = _RAND_2291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2292 = {1{`RANDOM}};
  _T_1334_re = _RAND_2292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2293 = {1{`RANDOM}};
  _T_1334_im = _RAND_2293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2294 = {1{`RANDOM}};
  _T_1335_re = _RAND_2294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2295 = {1{`RANDOM}};
  _T_1335_im = _RAND_2295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2296 = {1{`RANDOM}};
  _T_1336_re = _RAND_2296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2297 = {1{`RANDOM}};
  _T_1336_im = _RAND_2297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2298 = {1{`RANDOM}};
  _T_1337_re = _RAND_2298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2299 = {1{`RANDOM}};
  _T_1337_im = _RAND_2299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2300 = {1{`RANDOM}};
  _T_1338_re = _RAND_2300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2301 = {1{`RANDOM}};
  _T_1338_im = _RAND_2301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2302 = {1{`RANDOM}};
  _T_1339_re = _RAND_2302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2303 = {1{`RANDOM}};
  _T_1339_im = _RAND_2303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2304 = {1{`RANDOM}};
  _T_1340_re = _RAND_2304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2305 = {1{`RANDOM}};
  _T_1340_im = _RAND_2305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2306 = {1{`RANDOM}};
  _T_1341_re = _RAND_2306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2307 = {1{`RANDOM}};
  _T_1341_im = _RAND_2307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2308 = {1{`RANDOM}};
  _T_1342_re = _RAND_2308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2309 = {1{`RANDOM}};
  _T_1342_im = _RAND_2309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2310 = {1{`RANDOM}};
  _T_1343_re = _RAND_2310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2311 = {1{`RANDOM}};
  _T_1343_im = _RAND_2311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2312 = {1{`RANDOM}};
  _T_1344_re = _RAND_2312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2313 = {1{`RANDOM}};
  _T_1344_im = _RAND_2313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2314 = {1{`RANDOM}};
  _T_1345_re = _RAND_2314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2315 = {1{`RANDOM}};
  _T_1345_im = _RAND_2315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2316 = {1{`RANDOM}};
  _T_1346_re = _RAND_2316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2317 = {1{`RANDOM}};
  _T_1346_im = _RAND_2317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2318 = {1{`RANDOM}};
  _T_1347_re = _RAND_2318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2319 = {1{`RANDOM}};
  _T_1347_im = _RAND_2319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2320 = {1{`RANDOM}};
  _T_1348_re = _RAND_2320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2321 = {1{`RANDOM}};
  _T_1348_im = _RAND_2321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2322 = {1{`RANDOM}};
  _T_1349_re = _RAND_2322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2323 = {1{`RANDOM}};
  _T_1349_im = _RAND_2323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2324 = {1{`RANDOM}};
  _T_1350_re = _RAND_2324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2325 = {1{`RANDOM}};
  _T_1350_im = _RAND_2325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2326 = {1{`RANDOM}};
  _T_1351_re = _RAND_2326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2327 = {1{`RANDOM}};
  _T_1351_im = _RAND_2327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2328 = {1{`RANDOM}};
  _T_1352_re = _RAND_2328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2329 = {1{`RANDOM}};
  _T_1352_im = _RAND_2329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2330 = {1{`RANDOM}};
  _T_1353_re = _RAND_2330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2331 = {1{`RANDOM}};
  _T_1353_im = _RAND_2331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2332 = {1{`RANDOM}};
  _T_1354_re = _RAND_2332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2333 = {1{`RANDOM}};
  _T_1354_im = _RAND_2333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2334 = {1{`RANDOM}};
  _T_1355_re = _RAND_2334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2335 = {1{`RANDOM}};
  _T_1355_im = _RAND_2335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2336 = {1{`RANDOM}};
  _T_1356_re = _RAND_2336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2337 = {1{`RANDOM}};
  _T_1356_im = _RAND_2337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2338 = {1{`RANDOM}};
  _T_1357_re = _RAND_2338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2339 = {1{`RANDOM}};
  _T_1357_im = _RAND_2339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2340 = {1{`RANDOM}};
  _T_1358_re = _RAND_2340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2341 = {1{`RANDOM}};
  _T_1358_im = _RAND_2341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2342 = {1{`RANDOM}};
  _T_1359_re = _RAND_2342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2343 = {1{`RANDOM}};
  _T_1359_im = _RAND_2343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2344 = {1{`RANDOM}};
  _T_1360_re = _RAND_2344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2345 = {1{`RANDOM}};
  _T_1360_im = _RAND_2345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2346 = {1{`RANDOM}};
  _T_1361_re = _RAND_2346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2347 = {1{`RANDOM}};
  _T_1361_im = _RAND_2347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2348 = {1{`RANDOM}};
  _T_1362_re = _RAND_2348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2349 = {1{`RANDOM}};
  _T_1362_im = _RAND_2349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2350 = {1{`RANDOM}};
  _T_1363_re = _RAND_2350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2351 = {1{`RANDOM}};
  _T_1363_im = _RAND_2351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2352 = {1{`RANDOM}};
  _T_1364_re = _RAND_2352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2353 = {1{`RANDOM}};
  _T_1364_im = _RAND_2353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2354 = {1{`RANDOM}};
  _T_1365_re = _RAND_2354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2355 = {1{`RANDOM}};
  _T_1365_im = _RAND_2355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2356 = {1{`RANDOM}};
  _T_1366_re = _RAND_2356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2357 = {1{`RANDOM}};
  _T_1366_im = _RAND_2357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2358 = {1{`RANDOM}};
  _T_1367_re = _RAND_2358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2359 = {1{`RANDOM}};
  _T_1367_im = _RAND_2359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2360 = {1{`RANDOM}};
  _T_1368_re = _RAND_2360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2361 = {1{`RANDOM}};
  _T_1368_im = _RAND_2361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2362 = {1{`RANDOM}};
  _T_1369_re = _RAND_2362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2363 = {1{`RANDOM}};
  _T_1369_im = _RAND_2363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2364 = {1{`RANDOM}};
  _T_1370_re = _RAND_2364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2365 = {1{`RANDOM}};
  _T_1370_im = _RAND_2365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2366 = {1{`RANDOM}};
  _T_1371_re = _RAND_2366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2367 = {1{`RANDOM}};
  _T_1371_im = _RAND_2367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2368 = {1{`RANDOM}};
  _T_1372_re = _RAND_2368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2369 = {1{`RANDOM}};
  _T_1372_im = _RAND_2369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2370 = {1{`RANDOM}};
  _T_1373_re = _RAND_2370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2371 = {1{`RANDOM}};
  _T_1373_im = _RAND_2371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2372 = {1{`RANDOM}};
  _T_1374_re = _RAND_2372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2373 = {1{`RANDOM}};
  _T_1374_im = _RAND_2373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2374 = {1{`RANDOM}};
  _T_1375_re = _RAND_2374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2375 = {1{`RANDOM}};
  _T_1375_im = _RAND_2375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2376 = {1{`RANDOM}};
  _T_1376_re = _RAND_2376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2377 = {1{`RANDOM}};
  _T_1376_im = _RAND_2377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2378 = {1{`RANDOM}};
  _T_1377_re = _RAND_2378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2379 = {1{`RANDOM}};
  _T_1377_im = _RAND_2379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2380 = {1{`RANDOM}};
  _T_1378_re = _RAND_2380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2381 = {1{`RANDOM}};
  _T_1378_im = _RAND_2381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2382 = {1{`RANDOM}};
  _T_1379_re = _RAND_2382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2383 = {1{`RANDOM}};
  _T_1379_im = _RAND_2383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2384 = {1{`RANDOM}};
  _T_1380_re = _RAND_2384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2385 = {1{`RANDOM}};
  _T_1380_im = _RAND_2385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2386 = {1{`RANDOM}};
  _T_1381_re = _RAND_2386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2387 = {1{`RANDOM}};
  _T_1381_im = _RAND_2387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2388 = {1{`RANDOM}};
  _T_1382_re = _RAND_2388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2389 = {1{`RANDOM}};
  _T_1382_im = _RAND_2389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2390 = {1{`RANDOM}};
  _T_1383_re = _RAND_2390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2391 = {1{`RANDOM}};
  _T_1383_im = _RAND_2391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2392 = {1{`RANDOM}};
  _T_1384_re = _RAND_2392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2393 = {1{`RANDOM}};
  _T_1384_im = _RAND_2393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2394 = {1{`RANDOM}};
  _T_1385_re = _RAND_2394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2395 = {1{`RANDOM}};
  _T_1385_im = _RAND_2395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2396 = {1{`RANDOM}};
  _T_1386_re = _RAND_2396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2397 = {1{`RANDOM}};
  _T_1386_im = _RAND_2397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2398 = {1{`RANDOM}};
  _T_1387_re = _RAND_2398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2399 = {1{`RANDOM}};
  _T_1387_im = _RAND_2399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2400 = {1{`RANDOM}};
  _T_1388_re = _RAND_2400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2401 = {1{`RANDOM}};
  _T_1388_im = _RAND_2401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2402 = {1{`RANDOM}};
  _T_1389_re = _RAND_2402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2403 = {1{`RANDOM}};
  _T_1389_im = _RAND_2403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2404 = {1{`RANDOM}};
  _T_1390_re = _RAND_2404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2405 = {1{`RANDOM}};
  _T_1390_im = _RAND_2405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2406 = {1{`RANDOM}};
  _T_1391_re = _RAND_2406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2407 = {1{`RANDOM}};
  _T_1391_im = _RAND_2407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2408 = {1{`RANDOM}};
  _T_1392_re = _RAND_2408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2409 = {1{`RANDOM}};
  _T_1392_im = _RAND_2409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2410 = {1{`RANDOM}};
  _T_1393_re = _RAND_2410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2411 = {1{`RANDOM}};
  _T_1393_im = _RAND_2411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2412 = {1{`RANDOM}};
  _T_1394_re = _RAND_2412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2413 = {1{`RANDOM}};
  _T_1394_im = _RAND_2413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2414 = {1{`RANDOM}};
  _T_1395_re = _RAND_2414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2415 = {1{`RANDOM}};
  _T_1395_im = _RAND_2415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2416 = {1{`RANDOM}};
  _T_1396_re = _RAND_2416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2417 = {1{`RANDOM}};
  _T_1396_im = _RAND_2417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2418 = {1{`RANDOM}};
  _T_1397_re = _RAND_2418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2419 = {1{`RANDOM}};
  _T_1397_im = _RAND_2419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2420 = {1{`RANDOM}};
  _T_1398_re = _RAND_2420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2421 = {1{`RANDOM}};
  _T_1398_im = _RAND_2421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2422 = {1{`RANDOM}};
  _T_1399_re = _RAND_2422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2423 = {1{`RANDOM}};
  _T_1399_im = _RAND_2423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2424 = {1{`RANDOM}};
  _T_1400_re = _RAND_2424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2425 = {1{`RANDOM}};
  _T_1400_im = _RAND_2425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2426 = {1{`RANDOM}};
  _T_1401_re = _RAND_2426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2427 = {1{`RANDOM}};
  _T_1401_im = _RAND_2427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2428 = {1{`RANDOM}};
  _T_1402_re = _RAND_2428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2429 = {1{`RANDOM}};
  _T_1402_im = _RAND_2429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2430 = {1{`RANDOM}};
  _T_1403_re = _RAND_2430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2431 = {1{`RANDOM}};
  _T_1403_im = _RAND_2431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2432 = {1{`RANDOM}};
  _T_1404_re = _RAND_2432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2433 = {1{`RANDOM}};
  _T_1404_im = _RAND_2433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2434 = {1{`RANDOM}};
  _T_1405_re = _RAND_2434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2435 = {1{`RANDOM}};
  _T_1405_im = _RAND_2435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2436 = {1{`RANDOM}};
  _T_1406_re = _RAND_2436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2437 = {1{`RANDOM}};
  _T_1406_im = _RAND_2437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2438 = {1{`RANDOM}};
  _T_1407_re = _RAND_2438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2439 = {1{`RANDOM}};
  _T_1407_im = _RAND_2439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2440 = {1{`RANDOM}};
  _T_1408_re = _RAND_2440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2441 = {1{`RANDOM}};
  _T_1408_im = _RAND_2441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2442 = {1{`RANDOM}};
  _T_1409_re = _RAND_2442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2443 = {1{`RANDOM}};
  _T_1409_im = _RAND_2443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2444 = {1{`RANDOM}};
  _T_1410_re = _RAND_2444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2445 = {1{`RANDOM}};
  _T_1410_im = _RAND_2445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2446 = {1{`RANDOM}};
  _T_1411_re = _RAND_2446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2447 = {1{`RANDOM}};
  _T_1411_im = _RAND_2447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2448 = {1{`RANDOM}};
  _T_1412_re = _RAND_2448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2449 = {1{`RANDOM}};
  _T_1412_im = _RAND_2449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2450 = {1{`RANDOM}};
  _T_1413_re = _RAND_2450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2451 = {1{`RANDOM}};
  _T_1413_im = _RAND_2451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2452 = {1{`RANDOM}};
  _T_1414_re = _RAND_2452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2453 = {1{`RANDOM}};
  _T_1414_im = _RAND_2453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2454 = {1{`RANDOM}};
  _T_1415_re = _RAND_2454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2455 = {1{`RANDOM}};
  _T_1415_im = _RAND_2455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2456 = {1{`RANDOM}};
  _T_1416_re = _RAND_2456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2457 = {1{`RANDOM}};
  _T_1416_im = _RAND_2457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2458 = {1{`RANDOM}};
  _T_1417_re = _RAND_2458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2459 = {1{`RANDOM}};
  _T_1417_im = _RAND_2459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2460 = {1{`RANDOM}};
  _T_1418_re = _RAND_2460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2461 = {1{`RANDOM}};
  _T_1418_im = _RAND_2461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2462 = {1{`RANDOM}};
  _T_1419_re = _RAND_2462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2463 = {1{`RANDOM}};
  _T_1419_im = _RAND_2463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2464 = {1{`RANDOM}};
  _T_1420_re = _RAND_2464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2465 = {1{`RANDOM}};
  _T_1420_im = _RAND_2465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2466 = {1{`RANDOM}};
  _T_1421_re = _RAND_2466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2467 = {1{`RANDOM}};
  _T_1421_im = _RAND_2467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2468 = {1{`RANDOM}};
  _T_1422_re = _RAND_2468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2469 = {1{`RANDOM}};
  _T_1422_im = _RAND_2469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2470 = {1{`RANDOM}};
  _T_1423_re = _RAND_2470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2471 = {1{`RANDOM}};
  _T_1423_im = _RAND_2471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2472 = {1{`RANDOM}};
  _T_1424_re = _RAND_2472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2473 = {1{`RANDOM}};
  _T_1424_im = _RAND_2473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2474 = {1{`RANDOM}};
  _T_1425_re = _RAND_2474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2475 = {1{`RANDOM}};
  _T_1425_im = _RAND_2475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2476 = {1{`RANDOM}};
  _T_1426_re = _RAND_2476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2477 = {1{`RANDOM}};
  _T_1426_im = _RAND_2477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2478 = {1{`RANDOM}};
  _T_1427_re = _RAND_2478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2479 = {1{`RANDOM}};
  _T_1427_im = _RAND_2479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2480 = {1{`RANDOM}};
  _T_1428_re = _RAND_2480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2481 = {1{`RANDOM}};
  _T_1428_im = _RAND_2481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2482 = {1{`RANDOM}};
  _T_1429_re = _RAND_2482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2483 = {1{`RANDOM}};
  _T_1429_im = _RAND_2483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2484 = {1{`RANDOM}};
  _T_1430_re = _RAND_2484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2485 = {1{`RANDOM}};
  _T_1430_im = _RAND_2485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2486 = {1{`RANDOM}};
  _T_1431_re = _RAND_2486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2487 = {1{`RANDOM}};
  _T_1431_im = _RAND_2487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2488 = {1{`RANDOM}};
  _T_1432_re = _RAND_2488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2489 = {1{`RANDOM}};
  _T_1432_im = _RAND_2489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2490 = {1{`RANDOM}};
  _T_1433_re = _RAND_2490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2491 = {1{`RANDOM}};
  _T_1433_im = _RAND_2491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2492 = {1{`RANDOM}};
  _T_1434_re = _RAND_2492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2493 = {1{`RANDOM}};
  _T_1434_im = _RAND_2493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2494 = {1{`RANDOM}};
  _T_1435_re = _RAND_2494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2495 = {1{`RANDOM}};
  _T_1435_im = _RAND_2495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2496 = {1{`RANDOM}};
  _T_1436_re = _RAND_2496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2497 = {1{`RANDOM}};
  _T_1436_im = _RAND_2497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2498 = {1{`RANDOM}};
  _T_1437_re = _RAND_2498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2499 = {1{`RANDOM}};
  _T_1437_im = _RAND_2499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2500 = {1{`RANDOM}};
  _T_1438_re = _RAND_2500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2501 = {1{`RANDOM}};
  _T_1438_im = _RAND_2501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2502 = {1{`RANDOM}};
  _T_1439_re = _RAND_2502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2503 = {1{`RANDOM}};
  _T_1439_im = _RAND_2503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2504 = {1{`RANDOM}};
  _T_1440_re = _RAND_2504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2505 = {1{`RANDOM}};
  _T_1440_im = _RAND_2505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2506 = {1{`RANDOM}};
  _T_1441_re = _RAND_2506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2507 = {1{`RANDOM}};
  _T_1441_im = _RAND_2507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2508 = {1{`RANDOM}};
  _T_1442_re = _RAND_2508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2509 = {1{`RANDOM}};
  _T_1442_im = _RAND_2509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2510 = {1{`RANDOM}};
  _T_1443_re = _RAND_2510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2511 = {1{`RANDOM}};
  _T_1443_im = _RAND_2511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2512 = {1{`RANDOM}};
  _T_1444_re = _RAND_2512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2513 = {1{`RANDOM}};
  _T_1444_im = _RAND_2513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2514 = {1{`RANDOM}};
  _T_1445_re = _RAND_2514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2515 = {1{`RANDOM}};
  _T_1445_im = _RAND_2515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2516 = {1{`RANDOM}};
  _T_1446_re = _RAND_2516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2517 = {1{`RANDOM}};
  _T_1446_im = _RAND_2517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2518 = {1{`RANDOM}};
  _T_1447_re = _RAND_2518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2519 = {1{`RANDOM}};
  _T_1447_im = _RAND_2519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2520 = {1{`RANDOM}};
  _T_1448_re = _RAND_2520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2521 = {1{`RANDOM}};
  _T_1448_im = _RAND_2521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2522 = {1{`RANDOM}};
  _T_1449_re = _RAND_2522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2523 = {1{`RANDOM}};
  _T_1449_im = _RAND_2523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2524 = {1{`RANDOM}};
  _T_1450_re = _RAND_2524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2525 = {1{`RANDOM}};
  _T_1450_im = _RAND_2525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2526 = {1{`RANDOM}};
  _T_1451_re = _RAND_2526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2527 = {1{`RANDOM}};
  _T_1451_im = _RAND_2527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2528 = {1{`RANDOM}};
  _T_1452_re = _RAND_2528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2529 = {1{`RANDOM}};
  _T_1452_im = _RAND_2529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2530 = {1{`RANDOM}};
  _T_1453_re = _RAND_2530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2531 = {1{`RANDOM}};
  _T_1453_im = _RAND_2531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2532 = {1{`RANDOM}};
  _T_1454_re = _RAND_2532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2533 = {1{`RANDOM}};
  _T_1454_im = _RAND_2533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2534 = {1{`RANDOM}};
  _T_1455_re = _RAND_2534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2535 = {1{`RANDOM}};
  _T_1455_im = _RAND_2535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2536 = {1{`RANDOM}};
  _T_1456_re = _RAND_2536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2537 = {1{`RANDOM}};
  _T_1456_im = _RAND_2537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2538 = {1{`RANDOM}};
  _T_1457_re = _RAND_2538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2539 = {1{`RANDOM}};
  _T_1457_im = _RAND_2539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2540 = {1{`RANDOM}};
  _T_1458_re = _RAND_2540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2541 = {1{`RANDOM}};
  _T_1458_im = _RAND_2541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2542 = {1{`RANDOM}};
  _T_1459_re = _RAND_2542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2543 = {1{`RANDOM}};
  _T_1459_im = _RAND_2543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2544 = {1{`RANDOM}};
  _T_1460_re = _RAND_2544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2545 = {1{`RANDOM}};
  _T_1460_im = _RAND_2545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2546 = {1{`RANDOM}};
  _T_1461_re = _RAND_2546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2547 = {1{`RANDOM}};
  _T_1461_im = _RAND_2547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2548 = {1{`RANDOM}};
  _T_1462_re = _RAND_2548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2549 = {1{`RANDOM}};
  _T_1462_im = _RAND_2549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2550 = {1{`RANDOM}};
  _T_1463_re = _RAND_2550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2551 = {1{`RANDOM}};
  _T_1463_im = _RAND_2551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2552 = {1{`RANDOM}};
  _T_1464_re = _RAND_2552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2553 = {1{`RANDOM}};
  _T_1464_im = _RAND_2553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2554 = {1{`RANDOM}};
  _T_1465_re = _RAND_2554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2555 = {1{`RANDOM}};
  _T_1465_im = _RAND_2555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2556 = {1{`RANDOM}};
  _T_1466_re = _RAND_2556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2557 = {1{`RANDOM}};
  _T_1466_im = _RAND_2557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2558 = {1{`RANDOM}};
  _T_1467_re = _RAND_2558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2559 = {1{`RANDOM}};
  _T_1467_im = _RAND_2559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2560 = {1{`RANDOM}};
  _T_1468_re = _RAND_2560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2561 = {1{`RANDOM}};
  _T_1468_im = _RAND_2561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2562 = {1{`RANDOM}};
  _T_1469_re = _RAND_2562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2563 = {1{`RANDOM}};
  _T_1469_im = _RAND_2563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2564 = {1{`RANDOM}};
  _T_1470_re = _RAND_2564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2565 = {1{`RANDOM}};
  _T_1470_im = _RAND_2565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2566 = {1{`RANDOM}};
  _T_1471_re = _RAND_2566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2567 = {1{`RANDOM}};
  _T_1471_im = _RAND_2567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2568 = {1{`RANDOM}};
  _T_1472_re = _RAND_2568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2569 = {1{`RANDOM}};
  _T_1472_im = _RAND_2569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2570 = {1{`RANDOM}};
  _T_1473_re = _RAND_2570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2571 = {1{`RANDOM}};
  _T_1473_im = _RAND_2571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2572 = {1{`RANDOM}};
  _T_1474_re = _RAND_2572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2573 = {1{`RANDOM}};
  _T_1474_im = _RAND_2573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2574 = {1{`RANDOM}};
  _T_1475_re = _RAND_2574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2575 = {1{`RANDOM}};
  _T_1475_im = _RAND_2575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2576 = {1{`RANDOM}};
  _T_1476_re = _RAND_2576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2577 = {1{`RANDOM}};
  _T_1476_im = _RAND_2577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2578 = {1{`RANDOM}};
  _T_1477_re = _RAND_2578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2579 = {1{`RANDOM}};
  _T_1477_im = _RAND_2579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2580 = {1{`RANDOM}};
  _T_1478_re = _RAND_2580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2581 = {1{`RANDOM}};
  _T_1478_im = _RAND_2581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2582 = {1{`RANDOM}};
  _T_1479_re = _RAND_2582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2583 = {1{`RANDOM}};
  _T_1479_im = _RAND_2583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2584 = {1{`RANDOM}};
  _T_1480_re = _RAND_2584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2585 = {1{`RANDOM}};
  _T_1480_im = _RAND_2585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2586 = {1{`RANDOM}};
  _T_1481_re = _RAND_2586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2587 = {1{`RANDOM}};
  _T_1481_im = _RAND_2587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2588 = {1{`RANDOM}};
  _T_1482_re = _RAND_2588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2589 = {1{`RANDOM}};
  _T_1482_im = _RAND_2589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2590 = {1{`RANDOM}};
  _T_1483_re = _RAND_2590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2591 = {1{`RANDOM}};
  _T_1483_im = _RAND_2591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2592 = {1{`RANDOM}};
  _T_1484_re = _RAND_2592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2593 = {1{`RANDOM}};
  _T_1484_im = _RAND_2593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2594 = {1{`RANDOM}};
  _T_1485_re = _RAND_2594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2595 = {1{`RANDOM}};
  _T_1485_im = _RAND_2595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2596 = {1{`RANDOM}};
  _T_1486_re = _RAND_2596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2597 = {1{`RANDOM}};
  _T_1486_im = _RAND_2597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2598 = {1{`RANDOM}};
  _T_1487_re = _RAND_2598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2599 = {1{`RANDOM}};
  _T_1487_im = _RAND_2599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2600 = {1{`RANDOM}};
  _T_1488_re = _RAND_2600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2601 = {1{`RANDOM}};
  _T_1488_im = _RAND_2601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2602 = {1{`RANDOM}};
  _T_1489_re = _RAND_2602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2603 = {1{`RANDOM}};
  _T_1489_im = _RAND_2603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2604 = {1{`RANDOM}};
  _T_1490_re = _RAND_2604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2605 = {1{`RANDOM}};
  _T_1490_im = _RAND_2605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2606 = {1{`RANDOM}};
  _T_1491_re = _RAND_2606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2607 = {1{`RANDOM}};
  _T_1491_im = _RAND_2607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2608 = {1{`RANDOM}};
  _T_1492_re = _RAND_2608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2609 = {1{`RANDOM}};
  _T_1492_im = _RAND_2609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2610 = {1{`RANDOM}};
  _T_1493_re = _RAND_2610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2611 = {1{`RANDOM}};
  _T_1493_im = _RAND_2611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2612 = {1{`RANDOM}};
  _T_1494_re = _RAND_2612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2613 = {1{`RANDOM}};
  _T_1494_im = _RAND_2613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2614 = {1{`RANDOM}};
  _T_1495_re = _RAND_2614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2615 = {1{`RANDOM}};
  _T_1495_im = _RAND_2615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2616 = {1{`RANDOM}};
  _T_1496_re = _RAND_2616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2617 = {1{`RANDOM}};
  _T_1496_im = _RAND_2617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2618 = {1{`RANDOM}};
  _T_1497_re = _RAND_2618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2619 = {1{`RANDOM}};
  _T_1497_im = _RAND_2619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2620 = {1{`RANDOM}};
  _T_1498_re = _RAND_2620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2621 = {1{`RANDOM}};
  _T_1498_im = _RAND_2621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2622 = {1{`RANDOM}};
  _T_1499_re = _RAND_2622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2623 = {1{`RANDOM}};
  _T_1499_im = _RAND_2623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2624 = {1{`RANDOM}};
  _T_1500_re = _RAND_2624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2625 = {1{`RANDOM}};
  _T_1500_im = _RAND_2625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2626 = {1{`RANDOM}};
  _T_1501_re = _RAND_2626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2627 = {1{`RANDOM}};
  _T_1501_im = _RAND_2627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2628 = {1{`RANDOM}};
  _T_1502_re = _RAND_2628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2629 = {1{`RANDOM}};
  _T_1502_im = _RAND_2629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2630 = {1{`RANDOM}};
  _T_1503_re = _RAND_2630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2631 = {1{`RANDOM}};
  _T_1503_im = _RAND_2631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2632 = {1{`RANDOM}};
  _T_1504_re = _RAND_2632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2633 = {1{`RANDOM}};
  _T_1504_im = _RAND_2633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2634 = {1{`RANDOM}};
  _T_1505_re = _RAND_2634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2635 = {1{`RANDOM}};
  _T_1505_im = _RAND_2635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2636 = {1{`RANDOM}};
  _T_1506_re = _RAND_2636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2637 = {1{`RANDOM}};
  _T_1506_im = _RAND_2637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2638 = {1{`RANDOM}};
  _T_1507_re = _RAND_2638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2639 = {1{`RANDOM}};
  _T_1507_im = _RAND_2639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2640 = {1{`RANDOM}};
  _T_1508_re = _RAND_2640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2641 = {1{`RANDOM}};
  _T_1508_im = _RAND_2641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2642 = {1{`RANDOM}};
  _T_1509_re = _RAND_2642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2643 = {1{`RANDOM}};
  _T_1509_im = _RAND_2643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2644 = {1{`RANDOM}};
  _T_1510_re = _RAND_2644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2645 = {1{`RANDOM}};
  _T_1510_im = _RAND_2645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2646 = {1{`RANDOM}};
  _T_1511_re = _RAND_2646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2647 = {1{`RANDOM}};
  _T_1511_im = _RAND_2647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2648 = {1{`RANDOM}};
  _T_1512_re = _RAND_2648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2649 = {1{`RANDOM}};
  _T_1512_im = _RAND_2649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2650 = {1{`RANDOM}};
  _T_1513_re = _RAND_2650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2651 = {1{`RANDOM}};
  _T_1513_im = _RAND_2651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2652 = {1{`RANDOM}};
  _T_1514_re = _RAND_2652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2653 = {1{`RANDOM}};
  _T_1514_im = _RAND_2653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2654 = {1{`RANDOM}};
  _T_1515_re = _RAND_2654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2655 = {1{`RANDOM}};
  _T_1515_im = _RAND_2655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2656 = {1{`RANDOM}};
  _T_1516_re = _RAND_2656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2657 = {1{`RANDOM}};
  _T_1516_im = _RAND_2657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2658 = {1{`RANDOM}};
  _T_1517_re = _RAND_2658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2659 = {1{`RANDOM}};
  _T_1517_im = _RAND_2659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2660 = {1{`RANDOM}};
  _T_1518_re = _RAND_2660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2661 = {1{`RANDOM}};
  _T_1518_im = _RAND_2661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2662 = {1{`RANDOM}};
  _T_1519_re = _RAND_2662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2663 = {1{`RANDOM}};
  _T_1519_im = _RAND_2663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2664 = {1{`RANDOM}};
  _T_1520_re = _RAND_2664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2665 = {1{`RANDOM}};
  _T_1520_im = _RAND_2665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2666 = {1{`RANDOM}};
  _T_1521_re = _RAND_2666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2667 = {1{`RANDOM}};
  _T_1521_im = _RAND_2667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2668 = {1{`RANDOM}};
  _T_1522_re = _RAND_2668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2669 = {1{`RANDOM}};
  _T_1522_im = _RAND_2669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2670 = {1{`RANDOM}};
  _T_1523_re = _RAND_2670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2671 = {1{`RANDOM}};
  _T_1523_im = _RAND_2671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2672 = {1{`RANDOM}};
  _T_1524_re = _RAND_2672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2673 = {1{`RANDOM}};
  _T_1524_im = _RAND_2673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2674 = {1{`RANDOM}};
  _T_1525_re = _RAND_2674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2675 = {1{`RANDOM}};
  _T_1525_im = _RAND_2675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2676 = {1{`RANDOM}};
  _T_1526_re = _RAND_2676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2677 = {1{`RANDOM}};
  _T_1526_im = _RAND_2677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2678 = {1{`RANDOM}};
  _T_1527_re = _RAND_2678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2679 = {1{`RANDOM}};
  _T_1527_im = _RAND_2679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2680 = {1{`RANDOM}};
  _T_1528_re = _RAND_2680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2681 = {1{`RANDOM}};
  _T_1528_im = _RAND_2681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2682 = {1{`RANDOM}};
  _T_1529_re = _RAND_2682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2683 = {1{`RANDOM}};
  _T_1529_im = _RAND_2683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2684 = {1{`RANDOM}};
  _T_1530_re = _RAND_2684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2685 = {1{`RANDOM}};
  _T_1530_im = _RAND_2685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2686 = {1{`RANDOM}};
  _T_1531_re = _RAND_2686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2687 = {1{`RANDOM}};
  _T_1531_im = _RAND_2687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2688 = {1{`RANDOM}};
  _T_1532_re = _RAND_2688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2689 = {1{`RANDOM}};
  _T_1532_im = _RAND_2689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2690 = {1{`RANDOM}};
  _T_1533_re = _RAND_2690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2691 = {1{`RANDOM}};
  _T_1533_im = _RAND_2691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2692 = {1{`RANDOM}};
  _T_1534_re = _RAND_2692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2693 = {1{`RANDOM}};
  _T_1534_im = _RAND_2693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2694 = {1{`RANDOM}};
  _T_1535_re = _RAND_2694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2695 = {1{`RANDOM}};
  _T_1535_im = _RAND_2695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2696 = {1{`RANDOM}};
  _T_1536_re = _RAND_2696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2697 = {1{`RANDOM}};
  _T_1536_im = _RAND_2697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2698 = {1{`RANDOM}};
  _T_1537_re = _RAND_2698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2699 = {1{`RANDOM}};
  _T_1537_im = _RAND_2699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2700 = {1{`RANDOM}};
  _T_1538_re = _RAND_2700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2701 = {1{`RANDOM}};
  _T_1538_im = _RAND_2701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2702 = {1{`RANDOM}};
  _T_1539_re = _RAND_2702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2703 = {1{`RANDOM}};
  _T_1539_im = _RAND_2703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2704 = {1{`RANDOM}};
  _T_1540_re = _RAND_2704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2705 = {1{`RANDOM}};
  _T_1540_im = _RAND_2705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2706 = {1{`RANDOM}};
  _T_1541_re = _RAND_2706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2707 = {1{`RANDOM}};
  _T_1541_im = _RAND_2707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2708 = {1{`RANDOM}};
  _T_1542_re = _RAND_2708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2709 = {1{`RANDOM}};
  _T_1542_im = _RAND_2709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2710 = {1{`RANDOM}};
  _T_1543_re = _RAND_2710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2711 = {1{`RANDOM}};
  _T_1543_im = _RAND_2711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2712 = {1{`RANDOM}};
  _T_1544_re = _RAND_2712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2713 = {1{`RANDOM}};
  _T_1544_im = _RAND_2713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2714 = {1{`RANDOM}};
  _T_1545_re = _RAND_2714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2715 = {1{`RANDOM}};
  _T_1545_im = _RAND_2715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2716 = {1{`RANDOM}};
  _T_1546_re = _RAND_2716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2717 = {1{`RANDOM}};
  _T_1546_im = _RAND_2717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2718 = {1{`RANDOM}};
  _T_1547_re = _RAND_2718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2719 = {1{`RANDOM}};
  _T_1547_im = _RAND_2719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2720 = {1{`RANDOM}};
  _T_1548_re = _RAND_2720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2721 = {1{`RANDOM}};
  _T_1548_im = _RAND_2721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2722 = {1{`RANDOM}};
  _T_1549_re = _RAND_2722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2723 = {1{`RANDOM}};
  _T_1549_im = _RAND_2723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2724 = {1{`RANDOM}};
  _T_1550_re = _RAND_2724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2725 = {1{`RANDOM}};
  _T_1550_im = _RAND_2725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2726 = {1{`RANDOM}};
  _T_1551_re = _RAND_2726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2727 = {1{`RANDOM}};
  _T_1551_im = _RAND_2727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2728 = {1{`RANDOM}};
  _T_1552_re = _RAND_2728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2729 = {1{`RANDOM}};
  _T_1552_im = _RAND_2729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2730 = {1{`RANDOM}};
  _T_1553_re = _RAND_2730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2731 = {1{`RANDOM}};
  _T_1553_im = _RAND_2731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2732 = {1{`RANDOM}};
  _T_1554_re = _RAND_2732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2733 = {1{`RANDOM}};
  _T_1554_im = _RAND_2733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2734 = {1{`RANDOM}};
  _T_1555_re = _RAND_2734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2735 = {1{`RANDOM}};
  _T_1555_im = _RAND_2735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2736 = {1{`RANDOM}};
  _T_1556_re = _RAND_2736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2737 = {1{`RANDOM}};
  _T_1556_im = _RAND_2737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2738 = {1{`RANDOM}};
  _T_1557_re = _RAND_2738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2739 = {1{`RANDOM}};
  _T_1557_im = _RAND_2739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2740 = {1{`RANDOM}};
  _T_1558_re = _RAND_2740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2741 = {1{`RANDOM}};
  _T_1558_im = _RAND_2741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2742 = {1{`RANDOM}};
  _T_1559_re = _RAND_2742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2743 = {1{`RANDOM}};
  _T_1559_im = _RAND_2743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2744 = {1{`RANDOM}};
  _T_1560_re = _RAND_2744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2745 = {1{`RANDOM}};
  _T_1560_im = _RAND_2745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2746 = {1{`RANDOM}};
  _T_1561_re = _RAND_2746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2747 = {1{`RANDOM}};
  _T_1561_im = _RAND_2747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2748 = {1{`RANDOM}};
  _T_1562_re = _RAND_2748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2749 = {1{`RANDOM}};
  _T_1562_im = _RAND_2749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2750 = {1{`RANDOM}};
  _T_1563_re = _RAND_2750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2751 = {1{`RANDOM}};
  _T_1563_im = _RAND_2751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2752 = {1{`RANDOM}};
  _T_1564_re = _RAND_2752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2753 = {1{`RANDOM}};
  _T_1564_im = _RAND_2753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2754 = {1{`RANDOM}};
  _T_1565_re = _RAND_2754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2755 = {1{`RANDOM}};
  _T_1565_im = _RAND_2755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2756 = {1{`RANDOM}};
  _T_1566_re = _RAND_2756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2757 = {1{`RANDOM}};
  _T_1566_im = _RAND_2757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2758 = {1{`RANDOM}};
  _T_1567_re = _RAND_2758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2759 = {1{`RANDOM}};
  _T_1567_im = _RAND_2759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2760 = {1{`RANDOM}};
  _T_1568_re = _RAND_2760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2761 = {1{`RANDOM}};
  _T_1568_im = _RAND_2761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2762 = {1{`RANDOM}};
  _T_1569_re = _RAND_2762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2763 = {1{`RANDOM}};
  _T_1569_im = _RAND_2763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2764 = {1{`RANDOM}};
  _T_1570_re = _RAND_2764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2765 = {1{`RANDOM}};
  _T_1570_im = _RAND_2765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2766 = {1{`RANDOM}};
  _T_1571_re = _RAND_2766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2767 = {1{`RANDOM}};
  _T_1571_im = _RAND_2767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2768 = {1{`RANDOM}};
  _T_1572_re = _RAND_2768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2769 = {1{`RANDOM}};
  _T_1572_im = _RAND_2769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2770 = {1{`RANDOM}};
  _T_1573_re = _RAND_2770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2771 = {1{`RANDOM}};
  _T_1573_im = _RAND_2771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2772 = {1{`RANDOM}};
  _T_1574_re = _RAND_2772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2773 = {1{`RANDOM}};
  _T_1574_im = _RAND_2773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2774 = {1{`RANDOM}};
  _T_1575_re = _RAND_2774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2775 = {1{`RANDOM}};
  _T_1575_im = _RAND_2775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2776 = {1{`RANDOM}};
  _T_1576_re = _RAND_2776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2777 = {1{`RANDOM}};
  _T_1576_im = _RAND_2777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2778 = {1{`RANDOM}};
  _T_1577_re = _RAND_2778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2779 = {1{`RANDOM}};
  _T_1577_im = _RAND_2779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2780 = {1{`RANDOM}};
  _T_1578_re = _RAND_2780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2781 = {1{`RANDOM}};
  _T_1578_im = _RAND_2781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2782 = {1{`RANDOM}};
  _T_1579_re = _RAND_2782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2783 = {1{`RANDOM}};
  _T_1579_im = _RAND_2783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2784 = {1{`RANDOM}};
  _T_1580_re = _RAND_2784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2785 = {1{`RANDOM}};
  _T_1580_im = _RAND_2785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2786 = {1{`RANDOM}};
  _T_1581_re = _RAND_2786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2787 = {1{`RANDOM}};
  _T_1581_im = _RAND_2787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2788 = {1{`RANDOM}};
  _T_1582_re = _RAND_2788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2789 = {1{`RANDOM}};
  _T_1582_im = _RAND_2789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2790 = {1{`RANDOM}};
  _T_1583_re = _RAND_2790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2791 = {1{`RANDOM}};
  _T_1583_im = _RAND_2791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2792 = {1{`RANDOM}};
  _T_1584_re = _RAND_2792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2793 = {1{`RANDOM}};
  _T_1584_im = _RAND_2793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2794 = {1{`RANDOM}};
  _T_1585_re = _RAND_2794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2795 = {1{`RANDOM}};
  _T_1585_im = _RAND_2795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2796 = {1{`RANDOM}};
  _T_1586_re = _RAND_2796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2797 = {1{`RANDOM}};
  _T_1586_im = _RAND_2797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2798 = {1{`RANDOM}};
  _T_1587_re = _RAND_2798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2799 = {1{`RANDOM}};
  _T_1587_im = _RAND_2799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2800 = {1{`RANDOM}};
  _T_1588_re = _RAND_2800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2801 = {1{`RANDOM}};
  _T_1588_im = _RAND_2801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2802 = {1{`RANDOM}};
  _T_1589_re = _RAND_2802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2803 = {1{`RANDOM}};
  _T_1589_im = _RAND_2803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2804 = {1{`RANDOM}};
  _T_1590_re = _RAND_2804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2805 = {1{`RANDOM}};
  _T_1590_im = _RAND_2805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2806 = {1{`RANDOM}};
  _T_1591_re = _RAND_2806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2807 = {1{`RANDOM}};
  _T_1591_im = _RAND_2807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2808 = {1{`RANDOM}};
  _T_1592_re = _RAND_2808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2809 = {1{`RANDOM}};
  _T_1592_im = _RAND_2809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2810 = {1{`RANDOM}};
  _T_1593_re = _RAND_2810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2811 = {1{`RANDOM}};
  _T_1593_im = _RAND_2811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2812 = {1{`RANDOM}};
  _T_1594_re = _RAND_2812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2813 = {1{`RANDOM}};
  _T_1594_im = _RAND_2813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2814 = {1{`RANDOM}};
  _T_1595_re = _RAND_2814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2815 = {1{`RANDOM}};
  _T_1595_im = _RAND_2815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2816 = {1{`RANDOM}};
  _T_1596_re = _RAND_2816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2817 = {1{`RANDOM}};
  _T_1596_im = _RAND_2817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2818 = {1{`RANDOM}};
  _T_1597_re = _RAND_2818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2819 = {1{`RANDOM}};
  _T_1597_im = _RAND_2819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2820 = {1{`RANDOM}};
  _T_1598_re = _RAND_2820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2821 = {1{`RANDOM}};
  _T_1598_im = _RAND_2821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2822 = {1{`RANDOM}};
  _T_1599_re = _RAND_2822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2823 = {1{`RANDOM}};
  _T_1599_im = _RAND_2823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2824 = {1{`RANDOM}};
  _T_1600_re = _RAND_2824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2825 = {1{`RANDOM}};
  _T_1600_im = _RAND_2825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2826 = {1{`RANDOM}};
  _T_1601_re = _RAND_2826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2827 = {1{`RANDOM}};
  _T_1601_im = _RAND_2827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2828 = {1{`RANDOM}};
  _T_1602_re = _RAND_2828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2829 = {1{`RANDOM}};
  _T_1602_im = _RAND_2829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2830 = {1{`RANDOM}};
  _T_1603_re = _RAND_2830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2831 = {1{`RANDOM}};
  _T_1603_im = _RAND_2831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2832 = {1{`RANDOM}};
  _T_1604_re = _RAND_2832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2833 = {1{`RANDOM}};
  _T_1604_im = _RAND_2833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2834 = {1{`RANDOM}};
  _T_1605_re = _RAND_2834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2835 = {1{`RANDOM}};
  _T_1605_im = _RAND_2835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2836 = {1{`RANDOM}};
  _T_1606_re = _RAND_2836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2837 = {1{`RANDOM}};
  _T_1606_im = _RAND_2837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2838 = {1{`RANDOM}};
  _T_1607_re = _RAND_2838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2839 = {1{`RANDOM}};
  _T_1607_im = _RAND_2839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2840 = {1{`RANDOM}};
  _T_1608_re = _RAND_2840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2841 = {1{`RANDOM}};
  _T_1608_im = _RAND_2841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2842 = {1{`RANDOM}};
  _T_1609_re = _RAND_2842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2843 = {1{`RANDOM}};
  _T_1609_im = _RAND_2843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2844 = {1{`RANDOM}};
  _T_1610_re = _RAND_2844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2845 = {1{`RANDOM}};
  _T_1610_im = _RAND_2845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2846 = {1{`RANDOM}};
  _T_1611_re = _RAND_2846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2847 = {1{`RANDOM}};
  _T_1611_im = _RAND_2847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2848 = {1{`RANDOM}};
  _T_1612_re = _RAND_2848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2849 = {1{`RANDOM}};
  _T_1612_im = _RAND_2849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2850 = {1{`RANDOM}};
  _T_1613_re = _RAND_2850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2851 = {1{`RANDOM}};
  _T_1613_im = _RAND_2851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2852 = {1{`RANDOM}};
  _T_1614_re = _RAND_2852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2853 = {1{`RANDOM}};
  _T_1614_im = _RAND_2853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2854 = {1{`RANDOM}};
  _T_1615_re = _RAND_2854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2855 = {1{`RANDOM}};
  _T_1615_im = _RAND_2855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2856 = {1{`RANDOM}};
  _T_1616_re = _RAND_2856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2857 = {1{`RANDOM}};
  _T_1616_im = _RAND_2857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2858 = {1{`RANDOM}};
  _T_1617_re = _RAND_2858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2859 = {1{`RANDOM}};
  _T_1617_im = _RAND_2859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2860 = {1{`RANDOM}};
  _T_1618_re = _RAND_2860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2861 = {1{`RANDOM}};
  _T_1618_im = _RAND_2861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2862 = {1{`RANDOM}};
  _T_1619_re = _RAND_2862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2863 = {1{`RANDOM}};
  _T_1619_im = _RAND_2863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2864 = {1{`RANDOM}};
  _T_1620_re = _RAND_2864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2865 = {1{`RANDOM}};
  _T_1620_im = _RAND_2865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2866 = {1{`RANDOM}};
  _T_1621_re = _RAND_2866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2867 = {1{`RANDOM}};
  _T_1621_im = _RAND_2867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2868 = {1{`RANDOM}};
  _T_1622_re = _RAND_2868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2869 = {1{`RANDOM}};
  _T_1622_im = _RAND_2869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2870 = {1{`RANDOM}};
  _T_1623_re = _RAND_2870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2871 = {1{`RANDOM}};
  _T_1623_im = _RAND_2871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2872 = {1{`RANDOM}};
  _T_1624_re = _RAND_2872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2873 = {1{`RANDOM}};
  _T_1624_im = _RAND_2873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2874 = {1{`RANDOM}};
  _T_1625_re = _RAND_2874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2875 = {1{`RANDOM}};
  _T_1625_im = _RAND_2875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2876 = {1{`RANDOM}};
  _T_1626_re = _RAND_2876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2877 = {1{`RANDOM}};
  _T_1626_im = _RAND_2877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2878 = {1{`RANDOM}};
  _T_1627_re = _RAND_2878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2879 = {1{`RANDOM}};
  _T_1627_im = _RAND_2879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2880 = {1{`RANDOM}};
  _T_1628_re = _RAND_2880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2881 = {1{`RANDOM}};
  _T_1628_im = _RAND_2881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2882 = {1{`RANDOM}};
  _T_1629_re = _RAND_2882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2883 = {1{`RANDOM}};
  _T_1629_im = _RAND_2883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2884 = {1{`RANDOM}};
  _T_1630_re = _RAND_2884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2885 = {1{`RANDOM}};
  _T_1630_im = _RAND_2885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2886 = {1{`RANDOM}};
  _T_1631_re = _RAND_2886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2887 = {1{`RANDOM}};
  _T_1631_im = _RAND_2887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2888 = {1{`RANDOM}};
  _T_1632_re = _RAND_2888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2889 = {1{`RANDOM}};
  _T_1632_im = _RAND_2889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2890 = {1{`RANDOM}};
  _T_1633_re = _RAND_2890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2891 = {1{`RANDOM}};
  _T_1633_im = _RAND_2891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2892 = {1{`RANDOM}};
  _T_1634_re = _RAND_2892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2893 = {1{`RANDOM}};
  _T_1634_im = _RAND_2893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2894 = {1{`RANDOM}};
  _T_1635_re = _RAND_2894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2895 = {1{`RANDOM}};
  _T_1635_im = _RAND_2895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2896 = {1{`RANDOM}};
  _T_1636_re = _RAND_2896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2897 = {1{`RANDOM}};
  _T_1636_im = _RAND_2897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2898 = {1{`RANDOM}};
  _T_1637_re = _RAND_2898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2899 = {1{`RANDOM}};
  _T_1637_im = _RAND_2899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2900 = {1{`RANDOM}};
  _T_1638_re = _RAND_2900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2901 = {1{`RANDOM}};
  _T_1638_im = _RAND_2901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2902 = {1{`RANDOM}};
  _T_1639_re = _RAND_2902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2903 = {1{`RANDOM}};
  _T_1639_im = _RAND_2903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2904 = {1{`RANDOM}};
  _T_1640_re = _RAND_2904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2905 = {1{`RANDOM}};
  _T_1640_im = _RAND_2905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2906 = {1{`RANDOM}};
  _T_1641_re = _RAND_2906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2907 = {1{`RANDOM}};
  _T_1641_im = _RAND_2907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2908 = {1{`RANDOM}};
  _T_1642_re = _RAND_2908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2909 = {1{`RANDOM}};
  _T_1642_im = _RAND_2909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2910 = {1{`RANDOM}};
  _T_1643_re = _RAND_2910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2911 = {1{`RANDOM}};
  _T_1643_im = _RAND_2911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2912 = {1{`RANDOM}};
  _T_1644_re = _RAND_2912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2913 = {1{`RANDOM}};
  _T_1644_im = _RAND_2913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2914 = {1{`RANDOM}};
  _T_1645_re = _RAND_2914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2915 = {1{`RANDOM}};
  _T_1645_im = _RAND_2915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2916 = {1{`RANDOM}};
  _T_1646_re = _RAND_2916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2917 = {1{`RANDOM}};
  _T_1646_im = _RAND_2917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2918 = {1{`RANDOM}};
  _T_1647_re = _RAND_2918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2919 = {1{`RANDOM}};
  _T_1647_im = _RAND_2919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2920 = {1{`RANDOM}};
  _T_1648_re = _RAND_2920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2921 = {1{`RANDOM}};
  _T_1648_im = _RAND_2921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2922 = {1{`RANDOM}};
  _T_1649_re = _RAND_2922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2923 = {1{`RANDOM}};
  _T_1649_im = _RAND_2923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2924 = {1{`RANDOM}};
  _T_1650_re = _RAND_2924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2925 = {1{`RANDOM}};
  _T_1650_im = _RAND_2925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2926 = {1{`RANDOM}};
  _T_1651_re = _RAND_2926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2927 = {1{`RANDOM}};
  _T_1651_im = _RAND_2927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2928 = {1{`RANDOM}};
  _T_1652_re = _RAND_2928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2929 = {1{`RANDOM}};
  _T_1652_im = _RAND_2929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2930 = {1{`RANDOM}};
  _T_1653_re = _RAND_2930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2931 = {1{`RANDOM}};
  _T_1653_im = _RAND_2931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2932 = {1{`RANDOM}};
  _T_1654_re = _RAND_2932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2933 = {1{`RANDOM}};
  _T_1654_im = _RAND_2933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2934 = {1{`RANDOM}};
  _T_1655_re = _RAND_2934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2935 = {1{`RANDOM}};
  _T_1655_im = _RAND_2935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2936 = {1{`RANDOM}};
  _T_1656_re = _RAND_2936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2937 = {1{`RANDOM}};
  _T_1656_im = _RAND_2937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2938 = {1{`RANDOM}};
  _T_1657_re = _RAND_2938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2939 = {1{`RANDOM}};
  _T_1657_im = _RAND_2939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2940 = {1{`RANDOM}};
  _T_1658_re = _RAND_2940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2941 = {1{`RANDOM}};
  _T_1658_im = _RAND_2941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2942 = {1{`RANDOM}};
  _T_1659_re = _RAND_2942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2943 = {1{`RANDOM}};
  _T_1659_im = _RAND_2943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2944 = {1{`RANDOM}};
  _T_1660_re = _RAND_2944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2945 = {1{`RANDOM}};
  _T_1660_im = _RAND_2945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2946 = {1{`RANDOM}};
  _T_1661_re = _RAND_2946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2947 = {1{`RANDOM}};
  _T_1661_im = _RAND_2947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2948 = {1{`RANDOM}};
  _T_1662_re = _RAND_2948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2949 = {1{`RANDOM}};
  _T_1662_im = _RAND_2949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2950 = {1{`RANDOM}};
  _T_1663_re = _RAND_2950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2951 = {1{`RANDOM}};
  _T_1663_im = _RAND_2951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2952 = {1{`RANDOM}};
  _T_1664_re = _RAND_2952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2953 = {1{`RANDOM}};
  _T_1664_im = _RAND_2953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2954 = {1{`RANDOM}};
  _T_1665_re = _RAND_2954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2955 = {1{`RANDOM}};
  _T_1665_im = _RAND_2955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2956 = {1{`RANDOM}};
  _T_1666_re = _RAND_2956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2957 = {1{`RANDOM}};
  _T_1666_im = _RAND_2957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2958 = {1{`RANDOM}};
  _T_1667_re = _RAND_2958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2959 = {1{`RANDOM}};
  _T_1667_im = _RAND_2959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2960 = {1{`RANDOM}};
  _T_1668_re = _RAND_2960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2961 = {1{`RANDOM}};
  _T_1668_im = _RAND_2961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2962 = {1{`RANDOM}};
  _T_1669_re = _RAND_2962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2963 = {1{`RANDOM}};
  _T_1669_im = _RAND_2963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2964 = {1{`RANDOM}};
  _T_1670_re = _RAND_2964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2965 = {1{`RANDOM}};
  _T_1670_im = _RAND_2965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2966 = {1{`RANDOM}};
  _T_1671_re = _RAND_2966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2967 = {1{`RANDOM}};
  _T_1671_im = _RAND_2967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2968 = {1{`RANDOM}};
  _T_1672_re = _RAND_2968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2969 = {1{`RANDOM}};
  _T_1672_im = _RAND_2969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2970 = {1{`RANDOM}};
  _T_1673_re = _RAND_2970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2971 = {1{`RANDOM}};
  _T_1673_im = _RAND_2971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2972 = {1{`RANDOM}};
  _T_1674_re = _RAND_2972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2973 = {1{`RANDOM}};
  _T_1674_im = _RAND_2973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2974 = {1{`RANDOM}};
  _T_1675_re = _RAND_2974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2975 = {1{`RANDOM}};
  _T_1675_im = _RAND_2975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2976 = {1{`RANDOM}};
  _T_1676_re = _RAND_2976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2977 = {1{`RANDOM}};
  _T_1676_im = _RAND_2977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2978 = {1{`RANDOM}};
  _T_1677_re = _RAND_2978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2979 = {1{`RANDOM}};
  _T_1677_im = _RAND_2979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2980 = {1{`RANDOM}};
  _T_1678_re = _RAND_2980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2981 = {1{`RANDOM}};
  _T_1678_im = _RAND_2981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2982 = {1{`RANDOM}};
  _T_1679_re = _RAND_2982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2983 = {1{`RANDOM}};
  _T_1679_im = _RAND_2983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2984 = {1{`RANDOM}};
  _T_1680_re = _RAND_2984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2985 = {1{`RANDOM}};
  _T_1680_im = _RAND_2985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2986 = {1{`RANDOM}};
  _T_1681_re = _RAND_2986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2987 = {1{`RANDOM}};
  _T_1681_im = _RAND_2987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2988 = {1{`RANDOM}};
  _T_1682_re = _RAND_2988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2989 = {1{`RANDOM}};
  _T_1682_im = _RAND_2989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2990 = {1{`RANDOM}};
  _T_1683_re = _RAND_2990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2991 = {1{`RANDOM}};
  _T_1683_im = _RAND_2991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2992 = {1{`RANDOM}};
  _T_1684_re = _RAND_2992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2993 = {1{`RANDOM}};
  _T_1684_im = _RAND_2993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2994 = {1{`RANDOM}};
  _T_1685_re = _RAND_2994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2995 = {1{`RANDOM}};
  _T_1685_im = _RAND_2995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2996 = {1{`RANDOM}};
  _T_1686_re = _RAND_2996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2997 = {1{`RANDOM}};
  _T_1686_im = _RAND_2997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2998 = {1{`RANDOM}};
  _T_1687_re = _RAND_2998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2999 = {1{`RANDOM}};
  _T_1687_im = _RAND_2999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3000 = {1{`RANDOM}};
  _T_1688_re = _RAND_3000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3001 = {1{`RANDOM}};
  _T_1688_im = _RAND_3001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3002 = {1{`RANDOM}};
  _T_1689_re = _RAND_3002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3003 = {1{`RANDOM}};
  _T_1689_im = _RAND_3003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3004 = {1{`RANDOM}};
  _T_1690_re = _RAND_3004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3005 = {1{`RANDOM}};
  _T_1690_im = _RAND_3005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3006 = {1{`RANDOM}};
  _T_1691_re = _RAND_3006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3007 = {1{`RANDOM}};
  _T_1691_im = _RAND_3007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3008 = {1{`RANDOM}};
  _T_1692_re = _RAND_3008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3009 = {1{`RANDOM}};
  _T_1692_im = _RAND_3009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3010 = {1{`RANDOM}};
  _T_1693_re = _RAND_3010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3011 = {1{`RANDOM}};
  _T_1693_im = _RAND_3011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3012 = {1{`RANDOM}};
  _T_1694_re = _RAND_3012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3013 = {1{`RANDOM}};
  _T_1694_im = _RAND_3013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3014 = {1{`RANDOM}};
  _T_1695_re = _RAND_3014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3015 = {1{`RANDOM}};
  _T_1695_im = _RAND_3015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3016 = {1{`RANDOM}};
  _T_1696_re = _RAND_3016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3017 = {1{`RANDOM}};
  _T_1696_im = _RAND_3017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3018 = {1{`RANDOM}};
  _T_1697_re = _RAND_3018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3019 = {1{`RANDOM}};
  _T_1697_im = _RAND_3019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3020 = {1{`RANDOM}};
  _T_1698_re = _RAND_3020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3021 = {1{`RANDOM}};
  _T_1698_im = _RAND_3021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3022 = {1{`RANDOM}};
  _T_1699_re = _RAND_3022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3023 = {1{`RANDOM}};
  _T_1699_im = _RAND_3023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3024 = {1{`RANDOM}};
  _T_1700_re = _RAND_3024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3025 = {1{`RANDOM}};
  _T_1700_im = _RAND_3025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3026 = {1{`RANDOM}};
  _T_1701_re = _RAND_3026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3027 = {1{`RANDOM}};
  _T_1701_im = _RAND_3027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3028 = {1{`RANDOM}};
  _T_1702_re = _RAND_3028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3029 = {1{`RANDOM}};
  _T_1702_im = _RAND_3029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3030 = {1{`RANDOM}};
  _T_1703_re = _RAND_3030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3031 = {1{`RANDOM}};
  _T_1703_im = _RAND_3031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3032 = {1{`RANDOM}};
  _T_1704_re = _RAND_3032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3033 = {1{`RANDOM}};
  _T_1704_im = _RAND_3033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3034 = {1{`RANDOM}};
  _T_1705_re = _RAND_3034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3035 = {1{`RANDOM}};
  _T_1705_im = _RAND_3035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3036 = {1{`RANDOM}};
  _T_1706_re = _RAND_3036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3037 = {1{`RANDOM}};
  _T_1706_im = _RAND_3037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3038 = {1{`RANDOM}};
  _T_1707_re = _RAND_3038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3039 = {1{`RANDOM}};
  _T_1707_im = _RAND_3039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3040 = {1{`RANDOM}};
  _T_1708_re = _RAND_3040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3041 = {1{`RANDOM}};
  _T_1708_im = _RAND_3041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3042 = {1{`RANDOM}};
  _T_1709_re = _RAND_3042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3043 = {1{`RANDOM}};
  _T_1709_im = _RAND_3043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3044 = {1{`RANDOM}};
  _T_1710_re = _RAND_3044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3045 = {1{`RANDOM}};
  _T_1710_im = _RAND_3045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3046 = {1{`RANDOM}};
  _T_1711_re = _RAND_3046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3047 = {1{`RANDOM}};
  _T_1711_im = _RAND_3047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3048 = {1{`RANDOM}};
  _T_1712_re = _RAND_3048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3049 = {1{`RANDOM}};
  _T_1712_im = _RAND_3049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3050 = {1{`RANDOM}};
  _T_1713_re = _RAND_3050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3051 = {1{`RANDOM}};
  _T_1713_im = _RAND_3051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3052 = {1{`RANDOM}};
  _T_1714_re = _RAND_3052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3053 = {1{`RANDOM}};
  _T_1714_im = _RAND_3053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3054 = {1{`RANDOM}};
  _T_1715_re = _RAND_3054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3055 = {1{`RANDOM}};
  _T_1715_im = _RAND_3055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3056 = {1{`RANDOM}};
  _T_1716_re = _RAND_3056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3057 = {1{`RANDOM}};
  _T_1716_im = _RAND_3057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3058 = {1{`RANDOM}};
  _T_1717_re = _RAND_3058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3059 = {1{`RANDOM}};
  _T_1717_im = _RAND_3059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3060 = {1{`RANDOM}};
  _T_1718_re = _RAND_3060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3061 = {1{`RANDOM}};
  _T_1718_im = _RAND_3061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3062 = {1{`RANDOM}};
  _T_1719_re = _RAND_3062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3063 = {1{`RANDOM}};
  _T_1719_im = _RAND_3063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3064 = {1{`RANDOM}};
  _T_1720_re = _RAND_3064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3065 = {1{`RANDOM}};
  _T_1720_im = _RAND_3065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3066 = {1{`RANDOM}};
  _T_1721_re = _RAND_3066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3067 = {1{`RANDOM}};
  _T_1721_im = _RAND_3067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3068 = {1{`RANDOM}};
  _T_1722_re = _RAND_3068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3069 = {1{`RANDOM}};
  _T_1722_im = _RAND_3069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3070 = {1{`RANDOM}};
  _T_1723_re = _RAND_3070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3071 = {1{`RANDOM}};
  _T_1723_im = _RAND_3071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3072 = {1{`RANDOM}};
  _T_1724_re = _RAND_3072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3073 = {1{`RANDOM}};
  _T_1724_im = _RAND_3073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3074 = {1{`RANDOM}};
  _T_1725_re = _RAND_3074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3075 = {1{`RANDOM}};
  _T_1725_im = _RAND_3075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3076 = {1{`RANDOM}};
  _T_1726_re = _RAND_3076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3077 = {1{`RANDOM}};
  _T_1726_im = _RAND_3077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3078 = {1{`RANDOM}};
  _T_1727_re = _RAND_3078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3079 = {1{`RANDOM}};
  _T_1727_im = _RAND_3079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3080 = {1{`RANDOM}};
  _T_1728_re = _RAND_3080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3081 = {1{`RANDOM}};
  _T_1728_im = _RAND_3081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3082 = {1{`RANDOM}};
  _T_1729_re = _RAND_3082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3083 = {1{`RANDOM}};
  _T_1729_im = _RAND_3083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3084 = {1{`RANDOM}};
  _T_1730_re = _RAND_3084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3085 = {1{`RANDOM}};
  _T_1730_im = _RAND_3085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3086 = {1{`RANDOM}};
  _T_1731_re = _RAND_3086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3087 = {1{`RANDOM}};
  _T_1731_im = _RAND_3087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3088 = {1{`RANDOM}};
  _T_1732_re = _RAND_3088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3089 = {1{`RANDOM}};
  _T_1732_im = _RAND_3089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3090 = {1{`RANDOM}};
  _T_1733_re = _RAND_3090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3091 = {1{`RANDOM}};
  _T_1733_im = _RAND_3091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3092 = {1{`RANDOM}};
  _T_1734_re = _RAND_3092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3093 = {1{`RANDOM}};
  _T_1734_im = _RAND_3093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3094 = {1{`RANDOM}};
  _T_1735_re = _RAND_3094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3095 = {1{`RANDOM}};
  _T_1735_im = _RAND_3095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3096 = {1{`RANDOM}};
  _T_1736_re = _RAND_3096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3097 = {1{`RANDOM}};
  _T_1736_im = _RAND_3097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3098 = {1{`RANDOM}};
  _T_1737_re = _RAND_3098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3099 = {1{`RANDOM}};
  _T_1737_im = _RAND_3099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3100 = {1{`RANDOM}};
  _T_1738_re = _RAND_3100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3101 = {1{`RANDOM}};
  _T_1738_im = _RAND_3101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3102 = {1{`RANDOM}};
  _T_1739_re = _RAND_3102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3103 = {1{`RANDOM}};
  _T_1739_im = _RAND_3103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3104 = {1{`RANDOM}};
  _T_1740_re = _RAND_3104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3105 = {1{`RANDOM}};
  _T_1740_im = _RAND_3105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3106 = {1{`RANDOM}};
  _T_1741_re = _RAND_3106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3107 = {1{`RANDOM}};
  _T_1741_im = _RAND_3107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3108 = {1{`RANDOM}};
  _T_1742_re = _RAND_3108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3109 = {1{`RANDOM}};
  _T_1742_im = _RAND_3109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3110 = {1{`RANDOM}};
  _T_1743_re = _RAND_3110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3111 = {1{`RANDOM}};
  _T_1743_im = _RAND_3111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3112 = {1{`RANDOM}};
  _T_1744_re = _RAND_3112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3113 = {1{`RANDOM}};
  _T_1744_im = _RAND_3113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3114 = {1{`RANDOM}};
  _T_1745_re = _RAND_3114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3115 = {1{`RANDOM}};
  _T_1745_im = _RAND_3115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3116 = {1{`RANDOM}};
  _T_1746_re = _RAND_3116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3117 = {1{`RANDOM}};
  _T_1746_im = _RAND_3117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3118 = {1{`RANDOM}};
  _T_1747_re = _RAND_3118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3119 = {1{`RANDOM}};
  _T_1747_im = _RAND_3119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3120 = {1{`RANDOM}};
  _T_1748_re = _RAND_3120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3121 = {1{`RANDOM}};
  _T_1748_im = _RAND_3121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3122 = {1{`RANDOM}};
  _T_1749_re = _RAND_3122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3123 = {1{`RANDOM}};
  _T_1749_im = _RAND_3123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3124 = {1{`RANDOM}};
  _T_1750_re = _RAND_3124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3125 = {1{`RANDOM}};
  _T_1750_im = _RAND_3125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3126 = {1{`RANDOM}};
  _T_1751_re = _RAND_3126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3127 = {1{`RANDOM}};
  _T_1751_im = _RAND_3127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3128 = {1{`RANDOM}};
  _T_1752_re = _RAND_3128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3129 = {1{`RANDOM}};
  _T_1752_im = _RAND_3129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3130 = {1{`RANDOM}};
  _T_1753_re = _RAND_3130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3131 = {1{`RANDOM}};
  _T_1753_im = _RAND_3131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3132 = {1{`RANDOM}};
  _T_1754_re = _RAND_3132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3133 = {1{`RANDOM}};
  _T_1754_im = _RAND_3133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3134 = {1{`RANDOM}};
  _T_1755_re = _RAND_3134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3135 = {1{`RANDOM}};
  _T_1755_im = _RAND_3135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3136 = {1{`RANDOM}};
  _T_1756_re = _RAND_3136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3137 = {1{`RANDOM}};
  _T_1756_im = _RAND_3137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3138 = {1{`RANDOM}};
  _T_1757_re = _RAND_3138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3139 = {1{`RANDOM}};
  _T_1757_im = _RAND_3139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3140 = {1{`RANDOM}};
  _T_1758_re = _RAND_3140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3141 = {1{`RANDOM}};
  _T_1758_im = _RAND_3141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3142 = {1{`RANDOM}};
  _T_1759_re = _RAND_3142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3143 = {1{`RANDOM}};
  _T_1759_im = _RAND_3143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3144 = {1{`RANDOM}};
  _T_1760_re = _RAND_3144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3145 = {1{`RANDOM}};
  _T_1760_im = _RAND_3145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3146 = {1{`RANDOM}};
  _T_1761_re = _RAND_3146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3147 = {1{`RANDOM}};
  _T_1761_im = _RAND_3147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3148 = {1{`RANDOM}};
  _T_1762_re = _RAND_3148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3149 = {1{`RANDOM}};
  _T_1762_im = _RAND_3149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3150 = {1{`RANDOM}};
  _T_1763_re = _RAND_3150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3151 = {1{`RANDOM}};
  _T_1763_im = _RAND_3151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3152 = {1{`RANDOM}};
  _T_1764_re = _RAND_3152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3153 = {1{`RANDOM}};
  _T_1764_im = _RAND_3153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3154 = {1{`RANDOM}};
  _T_1765_re = _RAND_3154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3155 = {1{`RANDOM}};
  _T_1765_im = _RAND_3155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3156 = {1{`RANDOM}};
  _T_1766_re = _RAND_3156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3157 = {1{`RANDOM}};
  _T_1766_im = _RAND_3157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3158 = {1{`RANDOM}};
  _T_1767_re = _RAND_3158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3159 = {1{`RANDOM}};
  _T_1767_im = _RAND_3159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3160 = {1{`RANDOM}};
  _T_1768_re = _RAND_3160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3161 = {1{`RANDOM}};
  _T_1768_im = _RAND_3161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3162 = {1{`RANDOM}};
  _T_1769_re = _RAND_3162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3163 = {1{`RANDOM}};
  _T_1769_im = _RAND_3163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3164 = {1{`RANDOM}};
  _T_1770_re = _RAND_3164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3165 = {1{`RANDOM}};
  _T_1770_im = _RAND_3165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3166 = {1{`RANDOM}};
  _T_1771_re = _RAND_3166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3167 = {1{`RANDOM}};
  _T_1771_im = _RAND_3167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3168 = {1{`RANDOM}};
  _T_1772_re = _RAND_3168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3169 = {1{`RANDOM}};
  _T_1772_im = _RAND_3169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3170 = {1{`RANDOM}};
  _T_1773_re = _RAND_3170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3171 = {1{`RANDOM}};
  _T_1773_im = _RAND_3171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3172 = {1{`RANDOM}};
  _T_1774_re = _RAND_3172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3173 = {1{`RANDOM}};
  _T_1774_im = _RAND_3173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3174 = {1{`RANDOM}};
  _T_1775_re = _RAND_3174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3175 = {1{`RANDOM}};
  _T_1775_im = _RAND_3175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3176 = {1{`RANDOM}};
  _T_1776_re = _RAND_3176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3177 = {1{`RANDOM}};
  _T_1776_im = _RAND_3177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3178 = {1{`RANDOM}};
  _T_1777_re = _RAND_3178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3179 = {1{`RANDOM}};
  _T_1777_im = _RAND_3179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3180 = {1{`RANDOM}};
  _T_1778_re = _RAND_3180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3181 = {1{`RANDOM}};
  _T_1778_im = _RAND_3181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3182 = {1{`RANDOM}};
  _T_1779_re = _RAND_3182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3183 = {1{`RANDOM}};
  _T_1779_im = _RAND_3183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3184 = {1{`RANDOM}};
  _T_1780_re = _RAND_3184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3185 = {1{`RANDOM}};
  _T_1780_im = _RAND_3185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3186 = {1{`RANDOM}};
  _T_1781_re = _RAND_3186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3187 = {1{`RANDOM}};
  _T_1781_im = _RAND_3187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3188 = {1{`RANDOM}};
  _T_1782_re = _RAND_3188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3189 = {1{`RANDOM}};
  _T_1782_im = _RAND_3189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3190 = {1{`RANDOM}};
  _T_1783_re = _RAND_3190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3191 = {1{`RANDOM}};
  _T_1783_im = _RAND_3191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3192 = {1{`RANDOM}};
  _T_1784_re = _RAND_3192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3193 = {1{`RANDOM}};
  _T_1784_im = _RAND_3193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3194 = {1{`RANDOM}};
  _T_1785_re = _RAND_3194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3195 = {1{`RANDOM}};
  _T_1785_im = _RAND_3195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3196 = {1{`RANDOM}};
  _T_1786_re = _RAND_3196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3197 = {1{`RANDOM}};
  _T_1786_im = _RAND_3197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3198 = {1{`RANDOM}};
  _T_1787_re = _RAND_3198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3199 = {1{`RANDOM}};
  _T_1787_im = _RAND_3199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3200 = {1{`RANDOM}};
  _T_1788_re = _RAND_3200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3201 = {1{`RANDOM}};
  _T_1788_im = _RAND_3201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3202 = {1{`RANDOM}};
  _T_1789_re = _RAND_3202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3203 = {1{`RANDOM}};
  _T_1789_im = _RAND_3203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3204 = {1{`RANDOM}};
  _T_1790_re = _RAND_3204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3205 = {1{`RANDOM}};
  _T_1790_im = _RAND_3205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3206 = {1{`RANDOM}};
  _T_1791_re = _RAND_3206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3207 = {1{`RANDOM}};
  _T_1791_im = _RAND_3207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3208 = {1{`RANDOM}};
  _T_1792_re = _RAND_3208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3209 = {1{`RANDOM}};
  _T_1792_im = _RAND_3209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3210 = {1{`RANDOM}};
  _T_1793_re = _RAND_3210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3211 = {1{`RANDOM}};
  _T_1793_im = _RAND_3211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3212 = {1{`RANDOM}};
  _T_1794_re = _RAND_3212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3213 = {1{`RANDOM}};
  _T_1794_im = _RAND_3213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3214 = {1{`RANDOM}};
  _T_1795_re = _RAND_3214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3215 = {1{`RANDOM}};
  _T_1795_im = _RAND_3215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3216 = {1{`RANDOM}};
  _T_1796_re = _RAND_3216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3217 = {1{`RANDOM}};
  _T_1796_im = _RAND_3217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3218 = {1{`RANDOM}};
  _T_1797_re = _RAND_3218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3219 = {1{`RANDOM}};
  _T_1797_im = _RAND_3219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3220 = {1{`RANDOM}};
  _T_1798_re = _RAND_3220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3221 = {1{`RANDOM}};
  _T_1798_im = _RAND_3221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3222 = {1{`RANDOM}};
  _T_1799_re = _RAND_3222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3223 = {1{`RANDOM}};
  _T_1799_im = _RAND_3223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3224 = {1{`RANDOM}};
  _T_1800_re = _RAND_3224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3225 = {1{`RANDOM}};
  _T_1800_im = _RAND_3225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3226 = {1{`RANDOM}};
  _T_1801_re = _RAND_3226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3227 = {1{`RANDOM}};
  _T_1801_im = _RAND_3227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3228 = {1{`RANDOM}};
  _T_1802_re = _RAND_3228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3229 = {1{`RANDOM}};
  _T_1802_im = _RAND_3229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3230 = {1{`RANDOM}};
  _T_1803_re = _RAND_3230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3231 = {1{`RANDOM}};
  _T_1803_im = _RAND_3231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3232 = {1{`RANDOM}};
  _T_1804_re = _RAND_3232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3233 = {1{`RANDOM}};
  _T_1804_im = _RAND_3233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3234 = {1{`RANDOM}};
  _T_1805_re = _RAND_3234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3235 = {1{`RANDOM}};
  _T_1805_im = _RAND_3235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3236 = {1{`RANDOM}};
  _T_1806_re = _RAND_3236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3237 = {1{`RANDOM}};
  _T_1806_im = _RAND_3237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3238 = {1{`RANDOM}};
  _T_1807_re = _RAND_3238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3239 = {1{`RANDOM}};
  _T_1807_im = _RAND_3239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3240 = {1{`RANDOM}};
  _T_1808_re = _RAND_3240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3241 = {1{`RANDOM}};
  _T_1808_im = _RAND_3241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3242 = {1{`RANDOM}};
  _T_1809_re = _RAND_3242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3243 = {1{`RANDOM}};
  _T_1809_im = _RAND_3243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3244 = {1{`RANDOM}};
  _T_1810_re = _RAND_3244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3245 = {1{`RANDOM}};
  _T_1810_im = _RAND_3245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3246 = {1{`RANDOM}};
  _T_1811_re = _RAND_3246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3247 = {1{`RANDOM}};
  _T_1811_im = _RAND_3247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3248 = {1{`RANDOM}};
  _T_1812_re = _RAND_3248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3249 = {1{`RANDOM}};
  _T_1812_im = _RAND_3249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3250 = {1{`RANDOM}};
  _T_1813_re = _RAND_3250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3251 = {1{`RANDOM}};
  _T_1813_im = _RAND_3251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3252 = {1{`RANDOM}};
  _T_1814_re = _RAND_3252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3253 = {1{`RANDOM}};
  _T_1814_im = _RAND_3253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3254 = {1{`RANDOM}};
  _T_1815_re = _RAND_3254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3255 = {1{`RANDOM}};
  _T_1815_im = _RAND_3255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3256 = {1{`RANDOM}};
  _T_1816_re = _RAND_3256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3257 = {1{`RANDOM}};
  _T_1816_im = _RAND_3257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3258 = {1{`RANDOM}};
  _T_1817_re = _RAND_3258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3259 = {1{`RANDOM}};
  _T_1817_im = _RAND_3259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3260 = {1{`RANDOM}};
  _T_1818_re = _RAND_3260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3261 = {1{`RANDOM}};
  _T_1818_im = _RAND_3261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3262 = {1{`RANDOM}};
  _T_1819_re = _RAND_3262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3263 = {1{`RANDOM}};
  _T_1819_im = _RAND_3263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3264 = {1{`RANDOM}};
  _T_1820_re = _RAND_3264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3265 = {1{`RANDOM}};
  _T_1820_im = _RAND_3265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3266 = {1{`RANDOM}};
  _T_1821_re = _RAND_3266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3267 = {1{`RANDOM}};
  _T_1821_im = _RAND_3267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3268 = {1{`RANDOM}};
  _T_1822_re = _RAND_3268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3269 = {1{`RANDOM}};
  _T_1822_im = _RAND_3269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3270 = {1{`RANDOM}};
  _T_1823_re = _RAND_3270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3271 = {1{`RANDOM}};
  _T_1823_im = _RAND_3271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3272 = {1{`RANDOM}};
  _T_1824_re = _RAND_3272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3273 = {1{`RANDOM}};
  _T_1824_im = _RAND_3273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3274 = {1{`RANDOM}};
  _T_1825_re = _RAND_3274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3275 = {1{`RANDOM}};
  _T_1825_im = _RAND_3275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3276 = {1{`RANDOM}};
  _T_1826_re = _RAND_3276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3277 = {1{`RANDOM}};
  _T_1826_im = _RAND_3277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3278 = {1{`RANDOM}};
  _T_1827_re = _RAND_3278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3279 = {1{`RANDOM}};
  _T_1827_im = _RAND_3279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3280 = {1{`RANDOM}};
  _T_1828_re = _RAND_3280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3281 = {1{`RANDOM}};
  _T_1828_im = _RAND_3281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3282 = {1{`RANDOM}};
  _T_1829_re = _RAND_3282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3283 = {1{`RANDOM}};
  _T_1829_im = _RAND_3283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3284 = {1{`RANDOM}};
  _T_1830_re = _RAND_3284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3285 = {1{`RANDOM}};
  _T_1830_im = _RAND_3285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3286 = {1{`RANDOM}};
  _T_1831_re = _RAND_3286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3287 = {1{`RANDOM}};
  _T_1831_im = _RAND_3287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3288 = {1{`RANDOM}};
  _T_1832_re = _RAND_3288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3289 = {1{`RANDOM}};
  _T_1832_im = _RAND_3289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3290 = {1{`RANDOM}};
  _T_1833_re = _RAND_3290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3291 = {1{`RANDOM}};
  _T_1833_im = _RAND_3291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3292 = {1{`RANDOM}};
  _T_1834_re = _RAND_3292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3293 = {1{`RANDOM}};
  _T_1834_im = _RAND_3293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3294 = {1{`RANDOM}};
  _T_1835_re = _RAND_3294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3295 = {1{`RANDOM}};
  _T_1835_im = _RAND_3295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3296 = {1{`RANDOM}};
  _T_1836_re = _RAND_3296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3297 = {1{`RANDOM}};
  _T_1836_im = _RAND_3297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3298 = {1{`RANDOM}};
  _T_1837_re = _RAND_3298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3299 = {1{`RANDOM}};
  _T_1837_im = _RAND_3299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3300 = {1{`RANDOM}};
  _T_1838_re = _RAND_3300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3301 = {1{`RANDOM}};
  _T_1838_im = _RAND_3301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3302 = {1{`RANDOM}};
  _T_1839_re = _RAND_3302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3303 = {1{`RANDOM}};
  _T_1839_im = _RAND_3303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3304 = {1{`RANDOM}};
  _T_1840_re = _RAND_3304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3305 = {1{`RANDOM}};
  _T_1840_im = _RAND_3305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3306 = {1{`RANDOM}};
  _T_1841_re = _RAND_3306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3307 = {1{`RANDOM}};
  _T_1841_im = _RAND_3307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3308 = {1{`RANDOM}};
  _T_1842_re = _RAND_3308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3309 = {1{`RANDOM}};
  _T_1842_im = _RAND_3309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3310 = {1{`RANDOM}};
  _T_1843_re = _RAND_3310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3311 = {1{`RANDOM}};
  _T_1843_im = _RAND_3311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3312 = {1{`RANDOM}};
  _T_1844_re = _RAND_3312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3313 = {1{`RANDOM}};
  _T_1844_im = _RAND_3313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3314 = {1{`RANDOM}};
  _T_1845_re = _RAND_3314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3315 = {1{`RANDOM}};
  _T_1845_im = _RAND_3315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3316 = {1{`RANDOM}};
  _T_1846_re = _RAND_3316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3317 = {1{`RANDOM}};
  _T_1846_im = _RAND_3317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3318 = {1{`RANDOM}};
  _T_1847_re = _RAND_3318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3319 = {1{`RANDOM}};
  _T_1847_im = _RAND_3319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3320 = {1{`RANDOM}};
  _T_1848_re = _RAND_3320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3321 = {1{`RANDOM}};
  _T_1848_im = _RAND_3321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3322 = {1{`RANDOM}};
  _T_1849_re = _RAND_3322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3323 = {1{`RANDOM}};
  _T_1849_im = _RAND_3323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3324 = {1{`RANDOM}};
  _T_1850_re = _RAND_3324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3325 = {1{`RANDOM}};
  _T_1850_im = _RAND_3325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3326 = {1{`RANDOM}};
  _T_1851_re = _RAND_3326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3327 = {1{`RANDOM}};
  _T_1851_im = _RAND_3327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3328 = {1{`RANDOM}};
  _T_1852_re = _RAND_3328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3329 = {1{`RANDOM}};
  _T_1852_im = _RAND_3329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3330 = {1{`RANDOM}};
  _T_1853_re = _RAND_3330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3331 = {1{`RANDOM}};
  _T_1853_im = _RAND_3331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3332 = {1{`RANDOM}};
  _T_1854_re = _RAND_3332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3333 = {1{`RANDOM}};
  _T_1854_im = _RAND_3333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3334 = {1{`RANDOM}};
  _T_1855_re = _RAND_3334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3335 = {1{`RANDOM}};
  _T_1855_im = _RAND_3335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3336 = {1{`RANDOM}};
  _T_1856_re = _RAND_3336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3337 = {1{`RANDOM}};
  _T_1856_im = _RAND_3337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3338 = {1{`RANDOM}};
  _T_1857_re = _RAND_3338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3339 = {1{`RANDOM}};
  _T_1857_im = _RAND_3339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3340 = {1{`RANDOM}};
  _T_1858_re = _RAND_3340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3341 = {1{`RANDOM}};
  _T_1858_im = _RAND_3341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3342 = {1{`RANDOM}};
  _T_1859_re = _RAND_3342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3343 = {1{`RANDOM}};
  _T_1859_im = _RAND_3343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3344 = {1{`RANDOM}};
  _T_1860_re = _RAND_3344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3345 = {1{`RANDOM}};
  _T_1860_im = _RAND_3345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3346 = {1{`RANDOM}};
  _T_1861_re = _RAND_3346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3347 = {1{`RANDOM}};
  _T_1861_im = _RAND_3347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3348 = {1{`RANDOM}};
  _T_1862_re = _RAND_3348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3349 = {1{`RANDOM}};
  _T_1862_im = _RAND_3349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3350 = {1{`RANDOM}};
  _T_1863_re = _RAND_3350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3351 = {1{`RANDOM}};
  _T_1863_im = _RAND_3351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3352 = {1{`RANDOM}};
  _T_1864_re = _RAND_3352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3353 = {1{`RANDOM}};
  _T_1864_im = _RAND_3353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3354 = {1{`RANDOM}};
  _T_1865_re = _RAND_3354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3355 = {1{`RANDOM}};
  _T_1865_im = _RAND_3355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3356 = {1{`RANDOM}};
  _T_1866_re = _RAND_3356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3357 = {1{`RANDOM}};
  _T_1866_im = _RAND_3357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3358 = {1{`RANDOM}};
  _T_1867_re = _RAND_3358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3359 = {1{`RANDOM}};
  _T_1867_im = _RAND_3359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3360 = {1{`RANDOM}};
  _T_1868_re = _RAND_3360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3361 = {1{`RANDOM}};
  _T_1868_im = _RAND_3361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3362 = {1{`RANDOM}};
  _T_1869_re = _RAND_3362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3363 = {1{`RANDOM}};
  _T_1869_im = _RAND_3363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3364 = {1{`RANDOM}};
  _T_1870_re = _RAND_3364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3365 = {1{`RANDOM}};
  _T_1870_im = _RAND_3365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3366 = {1{`RANDOM}};
  _T_1871_re = _RAND_3366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3367 = {1{`RANDOM}};
  _T_1871_im = _RAND_3367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3368 = {1{`RANDOM}};
  _T_1872_re = _RAND_3368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3369 = {1{`RANDOM}};
  _T_1872_im = _RAND_3369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3370 = {1{`RANDOM}};
  _T_1873_re = _RAND_3370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3371 = {1{`RANDOM}};
  _T_1873_im = _RAND_3371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3372 = {1{`RANDOM}};
  _T_1874_re = _RAND_3372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3373 = {1{`RANDOM}};
  _T_1874_im = _RAND_3373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3374 = {1{`RANDOM}};
  _T_1875_re = _RAND_3374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3375 = {1{`RANDOM}};
  _T_1875_im = _RAND_3375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3376 = {1{`RANDOM}};
  _T_1876_re = _RAND_3376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3377 = {1{`RANDOM}};
  _T_1876_im = _RAND_3377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3378 = {1{`RANDOM}};
  _T_1877_re = _RAND_3378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3379 = {1{`RANDOM}};
  _T_1877_im = _RAND_3379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3380 = {1{`RANDOM}};
  _T_1878_re = _RAND_3380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3381 = {1{`RANDOM}};
  _T_1878_im = _RAND_3381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3382 = {1{`RANDOM}};
  _T_1879_re = _RAND_3382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3383 = {1{`RANDOM}};
  _T_1879_im = _RAND_3383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3384 = {1{`RANDOM}};
  _T_1880_re = _RAND_3384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3385 = {1{`RANDOM}};
  _T_1880_im = _RAND_3385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3386 = {1{`RANDOM}};
  _T_1881_re = _RAND_3386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3387 = {1{`RANDOM}};
  _T_1881_im = _RAND_3387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3388 = {1{`RANDOM}};
  _T_1882_re = _RAND_3388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3389 = {1{`RANDOM}};
  _T_1882_im = _RAND_3389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3390 = {1{`RANDOM}};
  _T_1883_re = _RAND_3390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3391 = {1{`RANDOM}};
  _T_1883_im = _RAND_3391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3392 = {1{`RANDOM}};
  _T_1884_re = _RAND_3392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3393 = {1{`RANDOM}};
  _T_1884_im = _RAND_3393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3394 = {1{`RANDOM}};
  _T_1885_re = _RAND_3394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3395 = {1{`RANDOM}};
  _T_1885_im = _RAND_3395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3396 = {1{`RANDOM}};
  _T_1886_re = _RAND_3396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3397 = {1{`RANDOM}};
  _T_1886_im = _RAND_3397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3398 = {1{`RANDOM}};
  _T_1887_re = _RAND_3398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3399 = {1{`RANDOM}};
  _T_1887_im = _RAND_3399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3400 = {1{`RANDOM}};
  _T_1888_re = _RAND_3400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3401 = {1{`RANDOM}};
  _T_1888_im = _RAND_3401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3402 = {1{`RANDOM}};
  _T_1889_re = _RAND_3402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3403 = {1{`RANDOM}};
  _T_1889_im = _RAND_3403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3404 = {1{`RANDOM}};
  _T_1890_re = _RAND_3404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3405 = {1{`RANDOM}};
  _T_1890_im = _RAND_3405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3406 = {1{`RANDOM}};
  _T_1891_re = _RAND_3406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3407 = {1{`RANDOM}};
  _T_1891_im = _RAND_3407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3408 = {1{`RANDOM}};
  _T_1892_re = _RAND_3408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3409 = {1{`RANDOM}};
  _T_1892_im = _RAND_3409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3410 = {1{`RANDOM}};
  _T_1893_re = _RAND_3410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3411 = {1{`RANDOM}};
  _T_1893_im = _RAND_3411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3412 = {1{`RANDOM}};
  _T_1894_re = _RAND_3412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3413 = {1{`RANDOM}};
  _T_1894_im = _RAND_3413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3414 = {1{`RANDOM}};
  _T_1895_re = _RAND_3414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3415 = {1{`RANDOM}};
  _T_1895_im = _RAND_3415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3416 = {1{`RANDOM}};
  _T_1896_re = _RAND_3416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3417 = {1{`RANDOM}};
  _T_1896_im = _RAND_3417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3418 = {1{`RANDOM}};
  _T_1897_re = _RAND_3418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3419 = {1{`RANDOM}};
  _T_1897_im = _RAND_3419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3420 = {1{`RANDOM}};
  _T_1898_re = _RAND_3420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3421 = {1{`RANDOM}};
  _T_1898_im = _RAND_3421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3422 = {1{`RANDOM}};
  _T_1899_re = _RAND_3422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3423 = {1{`RANDOM}};
  _T_1899_im = _RAND_3423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3424 = {1{`RANDOM}};
  _T_1900_re = _RAND_3424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3425 = {1{`RANDOM}};
  _T_1900_im = _RAND_3425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3426 = {1{`RANDOM}};
  _T_1901_re = _RAND_3426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3427 = {1{`RANDOM}};
  _T_1901_im = _RAND_3427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3428 = {1{`RANDOM}};
  _T_1902_re = _RAND_3428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3429 = {1{`RANDOM}};
  _T_1902_im = _RAND_3429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3430 = {1{`RANDOM}};
  _T_1903_re = _RAND_3430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3431 = {1{`RANDOM}};
  _T_1903_im = _RAND_3431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3432 = {1{`RANDOM}};
  _T_1904_re = _RAND_3432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3433 = {1{`RANDOM}};
  _T_1904_im = _RAND_3433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3434 = {1{`RANDOM}};
  _T_1905_re = _RAND_3434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3435 = {1{`RANDOM}};
  _T_1905_im = _RAND_3435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3436 = {1{`RANDOM}};
  _T_1906_re = _RAND_3436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3437 = {1{`RANDOM}};
  _T_1906_im = _RAND_3437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3438 = {1{`RANDOM}};
  _T_1907_re = _RAND_3438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3439 = {1{`RANDOM}};
  _T_1907_im = _RAND_3439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3440 = {1{`RANDOM}};
  _T_1908_re = _RAND_3440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3441 = {1{`RANDOM}};
  _T_1908_im = _RAND_3441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3442 = {1{`RANDOM}};
  _T_1909_re = _RAND_3442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3443 = {1{`RANDOM}};
  _T_1909_im = _RAND_3443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3444 = {1{`RANDOM}};
  _T_1910_re = _RAND_3444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3445 = {1{`RANDOM}};
  _T_1910_im = _RAND_3445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3446 = {1{`RANDOM}};
  _T_1911_re = _RAND_3446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3447 = {1{`RANDOM}};
  _T_1911_im = _RAND_3447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3448 = {1{`RANDOM}};
  _T_1912_re = _RAND_3448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3449 = {1{`RANDOM}};
  _T_1912_im = _RAND_3449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3450 = {1{`RANDOM}};
  _T_1913_re = _RAND_3450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3451 = {1{`RANDOM}};
  _T_1913_im = _RAND_3451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3452 = {1{`RANDOM}};
  _T_1914_re = _RAND_3452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3453 = {1{`RANDOM}};
  _T_1914_im = _RAND_3453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3454 = {1{`RANDOM}};
  _T_1915_re = _RAND_3454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3455 = {1{`RANDOM}};
  _T_1915_im = _RAND_3455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3456 = {1{`RANDOM}};
  _T_1916_re = _RAND_3456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3457 = {1{`RANDOM}};
  _T_1916_im = _RAND_3457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3458 = {1{`RANDOM}};
  _T_1917_re = _RAND_3458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3459 = {1{`RANDOM}};
  _T_1917_im = _RAND_3459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3460 = {1{`RANDOM}};
  _T_1918_re = _RAND_3460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3461 = {1{`RANDOM}};
  _T_1918_im = _RAND_3461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3462 = {1{`RANDOM}};
  _T_1919_re = _RAND_3462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3463 = {1{`RANDOM}};
  _T_1919_im = _RAND_3463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3464 = {1{`RANDOM}};
  _T_1920_re = _RAND_3464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3465 = {1{`RANDOM}};
  _T_1920_im = _RAND_3465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3466 = {1{`RANDOM}};
  _T_1921_re = _RAND_3466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3467 = {1{`RANDOM}};
  _T_1921_im = _RAND_3467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3468 = {1{`RANDOM}};
  _T_1922_re = _RAND_3468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3469 = {1{`RANDOM}};
  _T_1922_im = _RAND_3469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3470 = {1{`RANDOM}};
  _T_1923_re = _RAND_3470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3471 = {1{`RANDOM}};
  _T_1923_im = _RAND_3471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3472 = {1{`RANDOM}};
  _T_1924_re = _RAND_3472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3473 = {1{`RANDOM}};
  _T_1924_im = _RAND_3473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3474 = {1{`RANDOM}};
  _T_1925_re = _RAND_3474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3475 = {1{`RANDOM}};
  _T_1925_im = _RAND_3475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3476 = {1{`RANDOM}};
  _T_1926_re = _RAND_3476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3477 = {1{`RANDOM}};
  _T_1926_im = _RAND_3477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3478 = {1{`RANDOM}};
  _T_1927_re = _RAND_3478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3479 = {1{`RANDOM}};
  _T_1927_im = _RAND_3479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3480 = {1{`RANDOM}};
  _T_1928_re = _RAND_3480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3481 = {1{`RANDOM}};
  _T_1928_im = _RAND_3481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3482 = {1{`RANDOM}};
  _T_1929_re = _RAND_3482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3483 = {1{`RANDOM}};
  _T_1929_im = _RAND_3483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3484 = {1{`RANDOM}};
  _T_1930_re = _RAND_3484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3485 = {1{`RANDOM}};
  _T_1930_im = _RAND_3485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3486 = {1{`RANDOM}};
  _T_1931_re = _RAND_3486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3487 = {1{`RANDOM}};
  _T_1931_im = _RAND_3487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3488 = {1{`RANDOM}};
  _T_1932_re = _RAND_3488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3489 = {1{`RANDOM}};
  _T_1932_im = _RAND_3489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3490 = {1{`RANDOM}};
  _T_1933_re = _RAND_3490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3491 = {1{`RANDOM}};
  _T_1933_im = _RAND_3491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3492 = {1{`RANDOM}};
  _T_1934_re = _RAND_3492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3493 = {1{`RANDOM}};
  _T_1934_im = _RAND_3493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3494 = {1{`RANDOM}};
  _T_1935_re = _RAND_3494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3495 = {1{`RANDOM}};
  _T_1935_im = _RAND_3495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3496 = {1{`RANDOM}};
  _T_1936_re = _RAND_3496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3497 = {1{`RANDOM}};
  _T_1936_im = _RAND_3497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3498 = {1{`RANDOM}};
  _T_1937_re = _RAND_3498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3499 = {1{`RANDOM}};
  _T_1937_im = _RAND_3499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3500 = {1{`RANDOM}};
  _T_1938_re = _RAND_3500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3501 = {1{`RANDOM}};
  _T_1938_im = _RAND_3501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3502 = {1{`RANDOM}};
  _T_1939_re = _RAND_3502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3503 = {1{`RANDOM}};
  _T_1939_im = _RAND_3503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3504 = {1{`RANDOM}};
  _T_1940_re = _RAND_3504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3505 = {1{`RANDOM}};
  _T_1940_im = _RAND_3505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3506 = {1{`RANDOM}};
  _T_1941_re = _RAND_3506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3507 = {1{`RANDOM}};
  _T_1941_im = _RAND_3507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3508 = {1{`RANDOM}};
  _T_1942_re = _RAND_3508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3509 = {1{`RANDOM}};
  _T_1942_im = _RAND_3509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3510 = {1{`RANDOM}};
  _T_1943_re = _RAND_3510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3511 = {1{`RANDOM}};
  _T_1943_im = _RAND_3511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3512 = {1{`RANDOM}};
  _T_1944_re = _RAND_3512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3513 = {1{`RANDOM}};
  _T_1944_im = _RAND_3513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3514 = {1{`RANDOM}};
  _T_1945_re = _RAND_3514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3515 = {1{`RANDOM}};
  _T_1945_im = _RAND_3515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3516 = {1{`RANDOM}};
  _T_1946_re = _RAND_3516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3517 = {1{`RANDOM}};
  _T_1946_im = _RAND_3517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3518 = {1{`RANDOM}};
  _T_1947_re = _RAND_3518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3519 = {1{`RANDOM}};
  _T_1947_im = _RAND_3519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3520 = {1{`RANDOM}};
  _T_1948_re = _RAND_3520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3521 = {1{`RANDOM}};
  _T_1948_im = _RAND_3521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3522 = {1{`RANDOM}};
  _T_1949_re = _RAND_3522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3523 = {1{`RANDOM}};
  _T_1949_im = _RAND_3523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3524 = {1{`RANDOM}};
  _T_1950_re = _RAND_3524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3525 = {1{`RANDOM}};
  _T_1950_im = _RAND_3525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3526 = {1{`RANDOM}};
  _T_1951_re = _RAND_3526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3527 = {1{`RANDOM}};
  _T_1951_im = _RAND_3527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3528 = {1{`RANDOM}};
  _T_1952_re = _RAND_3528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3529 = {1{`RANDOM}};
  _T_1952_im = _RAND_3529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3530 = {1{`RANDOM}};
  _T_1953_re = _RAND_3530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3531 = {1{`RANDOM}};
  _T_1953_im = _RAND_3531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3532 = {1{`RANDOM}};
  _T_1954_re = _RAND_3532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3533 = {1{`RANDOM}};
  _T_1954_im = _RAND_3533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3534 = {1{`RANDOM}};
  _T_1955_re = _RAND_3534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3535 = {1{`RANDOM}};
  _T_1955_im = _RAND_3535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3536 = {1{`RANDOM}};
  _T_1956_re = _RAND_3536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3537 = {1{`RANDOM}};
  _T_1956_im = _RAND_3537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3538 = {1{`RANDOM}};
  _T_1957_re = _RAND_3538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3539 = {1{`RANDOM}};
  _T_1957_im = _RAND_3539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3540 = {1{`RANDOM}};
  _T_1958_re = _RAND_3540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3541 = {1{`RANDOM}};
  _T_1958_im = _RAND_3541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3542 = {1{`RANDOM}};
  _T_1959_re = _RAND_3542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3543 = {1{`RANDOM}};
  _T_1959_im = _RAND_3543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3544 = {1{`RANDOM}};
  _T_1960_re = _RAND_3544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3545 = {1{`RANDOM}};
  _T_1960_im = _RAND_3545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3546 = {1{`RANDOM}};
  _T_1961_re = _RAND_3546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3547 = {1{`RANDOM}};
  _T_1961_im = _RAND_3547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3548 = {1{`RANDOM}};
  _T_1962_re = _RAND_3548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3549 = {1{`RANDOM}};
  _T_1962_im = _RAND_3549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3550 = {1{`RANDOM}};
  _T_1963_re = _RAND_3550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3551 = {1{`RANDOM}};
  _T_1963_im = _RAND_3551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3552 = {1{`RANDOM}};
  _T_1964_re = _RAND_3552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3553 = {1{`RANDOM}};
  _T_1964_im = _RAND_3553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3554 = {1{`RANDOM}};
  _T_1965_re = _RAND_3554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3555 = {1{`RANDOM}};
  _T_1965_im = _RAND_3555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3556 = {1{`RANDOM}};
  _T_1966_re = _RAND_3556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3557 = {1{`RANDOM}};
  _T_1966_im = _RAND_3557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3558 = {1{`RANDOM}};
  _T_1967_re = _RAND_3558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3559 = {1{`RANDOM}};
  _T_1967_im = _RAND_3559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3560 = {1{`RANDOM}};
  _T_1968_re = _RAND_3560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3561 = {1{`RANDOM}};
  _T_1968_im = _RAND_3561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3562 = {1{`RANDOM}};
  _T_1969_re = _RAND_3562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3563 = {1{`RANDOM}};
  _T_1969_im = _RAND_3563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3564 = {1{`RANDOM}};
  _T_1970_re = _RAND_3564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3565 = {1{`RANDOM}};
  _T_1970_im = _RAND_3565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3566 = {1{`RANDOM}};
  _T_1971_re = _RAND_3566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3567 = {1{`RANDOM}};
  _T_1971_im = _RAND_3567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3568 = {1{`RANDOM}};
  _T_1972_re = _RAND_3568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3569 = {1{`RANDOM}};
  _T_1972_im = _RAND_3569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3570 = {1{`RANDOM}};
  _T_1973_re = _RAND_3570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3571 = {1{`RANDOM}};
  _T_1973_im = _RAND_3571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3572 = {1{`RANDOM}};
  _T_1974_re = _RAND_3572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3573 = {1{`RANDOM}};
  _T_1974_im = _RAND_3573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3574 = {1{`RANDOM}};
  _T_1975_re = _RAND_3574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3575 = {1{`RANDOM}};
  _T_1975_im = _RAND_3575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3576 = {1{`RANDOM}};
  _T_1976_re = _RAND_3576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3577 = {1{`RANDOM}};
  _T_1976_im = _RAND_3577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3578 = {1{`RANDOM}};
  _T_1977_re = _RAND_3578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3579 = {1{`RANDOM}};
  _T_1977_im = _RAND_3579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3580 = {1{`RANDOM}};
  _T_1978_re = _RAND_3580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3581 = {1{`RANDOM}};
  _T_1978_im = _RAND_3581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3582 = {1{`RANDOM}};
  _T_1979_re = _RAND_3582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3583 = {1{`RANDOM}};
  _T_1979_im = _RAND_3583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3584 = {1{`RANDOM}};
  _T_1980_re = _RAND_3584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3585 = {1{`RANDOM}};
  _T_1980_im = _RAND_3585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3586 = {1{`RANDOM}};
  _T_1981_re = _RAND_3586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3587 = {1{`RANDOM}};
  _T_1981_im = _RAND_3587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3588 = {1{`RANDOM}};
  _T_1982_re = _RAND_3588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3589 = {1{`RANDOM}};
  _T_1982_im = _RAND_3589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3590 = {1{`RANDOM}};
  _T_1983_re = _RAND_3590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3591 = {1{`RANDOM}};
  _T_1983_im = _RAND_3591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3592 = {1{`RANDOM}};
  _T_1984_re = _RAND_3592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3593 = {1{`RANDOM}};
  _T_1984_im = _RAND_3593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3594 = {1{`RANDOM}};
  _T_1985_re = _RAND_3594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3595 = {1{`RANDOM}};
  _T_1985_im = _RAND_3595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3596 = {1{`RANDOM}};
  _T_1986_re = _RAND_3596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3597 = {1{`RANDOM}};
  _T_1986_im = _RAND_3597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3598 = {1{`RANDOM}};
  _T_1987_re = _RAND_3598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3599 = {1{`RANDOM}};
  _T_1987_im = _RAND_3599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3600 = {1{`RANDOM}};
  _T_1988_re = _RAND_3600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3601 = {1{`RANDOM}};
  _T_1988_im = _RAND_3601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3602 = {1{`RANDOM}};
  _T_1989_re = _RAND_3602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3603 = {1{`RANDOM}};
  _T_1989_im = _RAND_3603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3604 = {1{`RANDOM}};
  _T_1990_re = _RAND_3604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3605 = {1{`RANDOM}};
  _T_1990_im = _RAND_3605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3606 = {1{`RANDOM}};
  _T_1991_re = _RAND_3606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3607 = {1{`RANDOM}};
  _T_1991_im = _RAND_3607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3608 = {1{`RANDOM}};
  _T_1992_re = _RAND_3608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3609 = {1{`RANDOM}};
  _T_1992_im = _RAND_3609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3610 = {1{`RANDOM}};
  _T_1993_re = _RAND_3610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3611 = {1{`RANDOM}};
  _T_1993_im = _RAND_3611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3612 = {1{`RANDOM}};
  _T_1994_re = _RAND_3612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3613 = {1{`RANDOM}};
  _T_1994_im = _RAND_3613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3614 = {1{`RANDOM}};
  _T_1995_re = _RAND_3614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3615 = {1{`RANDOM}};
  _T_1995_im = _RAND_3615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3616 = {1{`RANDOM}};
  _T_1996_re = _RAND_3616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3617 = {1{`RANDOM}};
  _T_1996_im = _RAND_3617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3618 = {1{`RANDOM}};
  _T_1997_re = _RAND_3618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3619 = {1{`RANDOM}};
  _T_1997_im = _RAND_3619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3620 = {1{`RANDOM}};
  _T_1998_re = _RAND_3620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3621 = {1{`RANDOM}};
  _T_1998_im = _RAND_3621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3622 = {1{`RANDOM}};
  _T_1999_re = _RAND_3622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3623 = {1{`RANDOM}};
  _T_1999_im = _RAND_3623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3624 = {1{`RANDOM}};
  _T_2000_re = _RAND_3624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3625 = {1{`RANDOM}};
  _T_2000_im = _RAND_3625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3626 = {1{`RANDOM}};
  _T_2001_re = _RAND_3626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3627 = {1{`RANDOM}};
  _T_2001_im = _RAND_3627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3628 = {1{`RANDOM}};
  _T_2002_re = _RAND_3628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3629 = {1{`RANDOM}};
  _T_2002_im = _RAND_3629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3630 = {1{`RANDOM}};
  _T_2003_re = _RAND_3630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3631 = {1{`RANDOM}};
  _T_2003_im = _RAND_3631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3632 = {1{`RANDOM}};
  _T_2004_re = _RAND_3632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3633 = {1{`RANDOM}};
  _T_2004_im = _RAND_3633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3634 = {1{`RANDOM}};
  _T_2005_re = _RAND_3634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3635 = {1{`RANDOM}};
  _T_2005_im = _RAND_3635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3636 = {1{`RANDOM}};
  _T_2006_re = _RAND_3636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3637 = {1{`RANDOM}};
  _T_2006_im = _RAND_3637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3638 = {1{`RANDOM}};
  _T_2007_re = _RAND_3638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3639 = {1{`RANDOM}};
  _T_2007_im = _RAND_3639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3640 = {1{`RANDOM}};
  _T_2008_re = _RAND_3640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3641 = {1{`RANDOM}};
  _T_2008_im = _RAND_3641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3642 = {1{`RANDOM}};
  _T_2009_re = _RAND_3642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3643 = {1{`RANDOM}};
  _T_2009_im = _RAND_3643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3644 = {1{`RANDOM}};
  _T_2010_re = _RAND_3644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3645 = {1{`RANDOM}};
  _T_2010_im = _RAND_3645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3646 = {1{`RANDOM}};
  _T_2011_re = _RAND_3646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3647 = {1{`RANDOM}};
  _T_2011_im = _RAND_3647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3648 = {1{`RANDOM}};
  _T_2012_re = _RAND_3648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3649 = {1{`RANDOM}};
  _T_2012_im = _RAND_3649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3650 = {1{`RANDOM}};
  _T_2013_re = _RAND_3650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3651 = {1{`RANDOM}};
  _T_2013_im = _RAND_3651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3652 = {1{`RANDOM}};
  _T_2014_re = _RAND_3652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3653 = {1{`RANDOM}};
  _T_2014_im = _RAND_3653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3654 = {1{`RANDOM}};
  _T_2015_re = _RAND_3654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3655 = {1{`RANDOM}};
  _T_2015_im = _RAND_3655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3656 = {1{`RANDOM}};
  _T_2016_re = _RAND_3656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3657 = {1{`RANDOM}};
  _T_2016_im = _RAND_3657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3658 = {1{`RANDOM}};
  _T_2017_re = _RAND_3658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3659 = {1{`RANDOM}};
  _T_2017_im = _RAND_3659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3660 = {1{`RANDOM}};
  _T_2018_re = _RAND_3660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3661 = {1{`RANDOM}};
  _T_2018_im = _RAND_3661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3662 = {1{`RANDOM}};
  _T_2019_re = _RAND_3662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3663 = {1{`RANDOM}};
  _T_2019_im = _RAND_3663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3664 = {1{`RANDOM}};
  _T_2020_re = _RAND_3664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3665 = {1{`RANDOM}};
  _T_2020_im = _RAND_3665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3666 = {1{`RANDOM}};
  _T_2021_re = _RAND_3666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3667 = {1{`RANDOM}};
  _T_2021_im = _RAND_3667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3668 = {1{`RANDOM}};
  _T_2022_re = _RAND_3668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3669 = {1{`RANDOM}};
  _T_2022_im = _RAND_3669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3670 = {1{`RANDOM}};
  _T_2023_re = _RAND_3670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3671 = {1{`RANDOM}};
  _T_2023_im = _RAND_3671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3672 = {1{`RANDOM}};
  _T_2024_re = _RAND_3672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3673 = {1{`RANDOM}};
  _T_2024_im = _RAND_3673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3674 = {1{`RANDOM}};
  _T_2025_re = _RAND_3674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3675 = {1{`RANDOM}};
  _T_2025_im = _RAND_3675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3676 = {1{`RANDOM}};
  _T_2026_re = _RAND_3676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3677 = {1{`RANDOM}};
  _T_2026_im = _RAND_3677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3678 = {1{`RANDOM}};
  _T_2027_re = _RAND_3678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3679 = {1{`RANDOM}};
  _T_2027_im = _RAND_3679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3680 = {1{`RANDOM}};
  _T_2028_re = _RAND_3680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3681 = {1{`RANDOM}};
  _T_2028_im = _RAND_3681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3682 = {1{`RANDOM}};
  _T_2029_re = _RAND_3682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3683 = {1{`RANDOM}};
  _T_2029_im = _RAND_3683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3684 = {1{`RANDOM}};
  _T_2030_re = _RAND_3684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3685 = {1{`RANDOM}};
  _T_2030_im = _RAND_3685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3686 = {1{`RANDOM}};
  _T_2031_re = _RAND_3686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3687 = {1{`RANDOM}};
  _T_2031_im = _RAND_3687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3688 = {1{`RANDOM}};
  _T_2032_re = _RAND_3688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3689 = {1{`RANDOM}};
  _T_2032_im = _RAND_3689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3690 = {1{`RANDOM}};
  _T_2033_re = _RAND_3690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3691 = {1{`RANDOM}};
  _T_2033_im = _RAND_3691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3692 = {1{`RANDOM}};
  _T_2034_re = _RAND_3692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3693 = {1{`RANDOM}};
  _T_2034_im = _RAND_3693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3694 = {1{`RANDOM}};
  _T_2035_re = _RAND_3694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3695 = {1{`RANDOM}};
  _T_2035_im = _RAND_3695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3696 = {1{`RANDOM}};
  _T_2036_re = _RAND_3696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3697 = {1{`RANDOM}};
  _T_2036_im = _RAND_3697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3698 = {1{`RANDOM}};
  _T_2037_re = _RAND_3698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3699 = {1{`RANDOM}};
  _T_2037_im = _RAND_3699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3700 = {1{`RANDOM}};
  _T_2038_re = _RAND_3700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3701 = {1{`RANDOM}};
  _T_2038_im = _RAND_3701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3702 = {1{`RANDOM}};
  _T_2039_re = _RAND_3702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3703 = {1{`RANDOM}};
  _T_2039_im = _RAND_3703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3704 = {1{`RANDOM}};
  _T_2040_re = _RAND_3704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3705 = {1{`RANDOM}};
  _T_2040_im = _RAND_3705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3706 = {1{`RANDOM}};
  _T_2041_re = _RAND_3706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3707 = {1{`RANDOM}};
  _T_2041_im = _RAND_3707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3708 = {1{`RANDOM}};
  _T_2042_re = _RAND_3708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3709 = {1{`RANDOM}};
  _T_2042_im = _RAND_3709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3710 = {1{`RANDOM}};
  _T_2043_re = _RAND_3710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3711 = {1{`RANDOM}};
  _T_2043_im = _RAND_3711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3712 = {1{`RANDOM}};
  _T_2044_re = _RAND_3712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3713 = {1{`RANDOM}};
  _T_2044_im = _RAND_3713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3714 = {1{`RANDOM}};
  _T_2045_re = _RAND_3714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3715 = {1{`RANDOM}};
  _T_2045_im = _RAND_3715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3716 = {1{`RANDOM}};
  _T_2046_re = _RAND_3716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3717 = {1{`RANDOM}};
  _T_2046_im = _RAND_3717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3718 = {1{`RANDOM}};
  _T_2047_re = _RAND_3718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3719 = {1{`RANDOM}};
  _T_2047_im = _RAND_3719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3720 = {1{`RANDOM}};
  _T_2048_re = _RAND_3720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3721 = {1{`RANDOM}};
  _T_2048_im = _RAND_3721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3722 = {1{`RANDOM}};
  _T_2049_re = _RAND_3722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3723 = {1{`RANDOM}};
  _T_2049_im = _RAND_3723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3724 = {1{`RANDOM}};
  _T_2050_re = _RAND_3724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3725 = {1{`RANDOM}};
  _T_2050_im = _RAND_3725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3726 = {1{`RANDOM}};
  _T_2051_re = _RAND_3726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3727 = {1{`RANDOM}};
  _T_2051_im = _RAND_3727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3728 = {1{`RANDOM}};
  _T_2052_re = _RAND_3728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3729 = {1{`RANDOM}};
  _T_2052_im = _RAND_3729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3730 = {1{`RANDOM}};
  _T_2053_re = _RAND_3730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3731 = {1{`RANDOM}};
  _T_2053_im = _RAND_3731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3732 = {1{`RANDOM}};
  _T_2054_re = _RAND_3732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3733 = {1{`RANDOM}};
  _T_2054_im = _RAND_3733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3734 = {1{`RANDOM}};
  _T_2055_re = _RAND_3734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3735 = {1{`RANDOM}};
  _T_2055_im = _RAND_3735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3736 = {1{`RANDOM}};
  _T_2056_re = _RAND_3736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3737 = {1{`RANDOM}};
  _T_2056_im = _RAND_3737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3738 = {1{`RANDOM}};
  _T_2057_re = _RAND_3738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3739 = {1{`RANDOM}};
  _T_2057_im = _RAND_3739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3740 = {1{`RANDOM}};
  _T_2058_re = _RAND_3740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3741 = {1{`RANDOM}};
  _T_2058_im = _RAND_3741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3742 = {1{`RANDOM}};
  _T_2059_re = _RAND_3742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3743 = {1{`RANDOM}};
  _T_2059_im = _RAND_3743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3744 = {1{`RANDOM}};
  _T_2060_re = _RAND_3744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3745 = {1{`RANDOM}};
  _T_2060_im = _RAND_3745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3746 = {1{`RANDOM}};
  _T_2061_re = _RAND_3746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3747 = {1{`RANDOM}};
  _T_2061_im = _RAND_3747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3748 = {1{`RANDOM}};
  _T_2062_re = _RAND_3748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3749 = {1{`RANDOM}};
  _T_2062_im = _RAND_3749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3750 = {1{`RANDOM}};
  _T_2063_re = _RAND_3750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3751 = {1{`RANDOM}};
  _T_2063_im = _RAND_3751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3752 = {1{`RANDOM}};
  _T_2064_re = _RAND_3752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3753 = {1{`RANDOM}};
  _T_2064_im = _RAND_3753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3754 = {1{`RANDOM}};
  _T_2065_re = _RAND_3754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3755 = {1{`RANDOM}};
  _T_2065_im = _RAND_3755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3756 = {1{`RANDOM}};
  _T_2066_re = _RAND_3756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3757 = {1{`RANDOM}};
  _T_2066_im = _RAND_3757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3758 = {1{`RANDOM}};
  _T_2067_re = _RAND_3758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3759 = {1{`RANDOM}};
  _T_2067_im = _RAND_3759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3760 = {1{`RANDOM}};
  _T_2068_re = _RAND_3760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3761 = {1{`RANDOM}};
  _T_2068_im = _RAND_3761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3762 = {1{`RANDOM}};
  _T_2069_re = _RAND_3762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3763 = {1{`RANDOM}};
  _T_2069_im = _RAND_3763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3764 = {1{`RANDOM}};
  _T_2070_re = _RAND_3764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3765 = {1{`RANDOM}};
  _T_2070_im = _RAND_3765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3766 = {1{`RANDOM}};
  _T_2071_re = _RAND_3766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3767 = {1{`RANDOM}};
  _T_2071_im = _RAND_3767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3768 = {1{`RANDOM}};
  _T_2072_re = _RAND_3768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3769 = {1{`RANDOM}};
  _T_2072_im = _RAND_3769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3770 = {1{`RANDOM}};
  _T_2073_re = _RAND_3770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3771 = {1{`RANDOM}};
  _T_2073_im = _RAND_3771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3772 = {1{`RANDOM}};
  _T_2074_re = _RAND_3772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3773 = {1{`RANDOM}};
  _T_2074_im = _RAND_3773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3774 = {1{`RANDOM}};
  _T_2075_re = _RAND_3774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3775 = {1{`RANDOM}};
  _T_2075_im = _RAND_3775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3776 = {1{`RANDOM}};
  _T_2076_re = _RAND_3776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3777 = {1{`RANDOM}};
  _T_2076_im = _RAND_3777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3778 = {1{`RANDOM}};
  _T_2077_re = _RAND_3778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3779 = {1{`RANDOM}};
  _T_2077_im = _RAND_3779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3780 = {1{`RANDOM}};
  _T_2078_re = _RAND_3780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3781 = {1{`RANDOM}};
  _T_2078_im = _RAND_3781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3782 = {1{`RANDOM}};
  _T_2079_re = _RAND_3782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3783 = {1{`RANDOM}};
  _T_2079_im = _RAND_3783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3784 = {1{`RANDOM}};
  _T_2080_re = _RAND_3784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3785 = {1{`RANDOM}};
  _T_2080_im = _RAND_3785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3786 = {1{`RANDOM}};
  _T_2081_re = _RAND_3786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3787 = {1{`RANDOM}};
  _T_2081_im = _RAND_3787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3788 = {1{`RANDOM}};
  _T_2082_re = _RAND_3788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3789 = {1{`RANDOM}};
  _T_2082_im = _RAND_3789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3790 = {1{`RANDOM}};
  _T_2083_re = _RAND_3790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3791 = {1{`RANDOM}};
  _T_2083_im = _RAND_3791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3792 = {1{`RANDOM}};
  _T_2084_re = _RAND_3792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3793 = {1{`RANDOM}};
  _T_2084_im = _RAND_3793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3794 = {1{`RANDOM}};
  _T_2085_re = _RAND_3794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3795 = {1{`RANDOM}};
  _T_2085_im = _RAND_3795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3796 = {1{`RANDOM}};
  _T_2086_re = _RAND_3796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3797 = {1{`RANDOM}};
  _T_2086_im = _RAND_3797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3798 = {1{`RANDOM}};
  _T_2087_re = _RAND_3798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3799 = {1{`RANDOM}};
  _T_2087_im = _RAND_3799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3800 = {1{`RANDOM}};
  _T_2088_re = _RAND_3800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3801 = {1{`RANDOM}};
  _T_2088_im = _RAND_3801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3802 = {1{`RANDOM}};
  _T_2089_re = _RAND_3802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3803 = {1{`RANDOM}};
  _T_2089_im = _RAND_3803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3804 = {1{`RANDOM}};
  _T_2090_re = _RAND_3804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3805 = {1{`RANDOM}};
  _T_2090_im = _RAND_3805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3806 = {1{`RANDOM}};
  _T_2091_re = _RAND_3806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3807 = {1{`RANDOM}};
  _T_2091_im = _RAND_3807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3808 = {1{`RANDOM}};
  _T_2092_re = _RAND_3808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3809 = {1{`RANDOM}};
  _T_2092_im = _RAND_3809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3810 = {1{`RANDOM}};
  _T_2093_re = _RAND_3810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3811 = {1{`RANDOM}};
  _T_2093_im = _RAND_3811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3812 = {1{`RANDOM}};
  _T_2094_re = _RAND_3812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3813 = {1{`RANDOM}};
  _T_2094_im = _RAND_3813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3814 = {1{`RANDOM}};
  _T_2095_re = _RAND_3814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3815 = {1{`RANDOM}};
  _T_2095_im = _RAND_3815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3816 = {1{`RANDOM}};
  _T_2096_re = _RAND_3816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3817 = {1{`RANDOM}};
  _T_2096_im = _RAND_3817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3818 = {1{`RANDOM}};
  _T_2097_re = _RAND_3818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3819 = {1{`RANDOM}};
  _T_2097_im = _RAND_3819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3820 = {1{`RANDOM}};
  _T_2098_re = _RAND_3820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3821 = {1{`RANDOM}};
  _T_2098_im = _RAND_3821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3822 = {1{`RANDOM}};
  _T_2099_re = _RAND_3822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3823 = {1{`RANDOM}};
  _T_2099_im = _RAND_3823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3824 = {1{`RANDOM}};
  _T_2100_re = _RAND_3824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3825 = {1{`RANDOM}};
  _T_2100_im = _RAND_3825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3826 = {1{`RANDOM}};
  _T_2101_re = _RAND_3826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3827 = {1{`RANDOM}};
  _T_2101_im = _RAND_3827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3828 = {1{`RANDOM}};
  _T_2102_re = _RAND_3828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3829 = {1{`RANDOM}};
  _T_2102_im = _RAND_3829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3830 = {1{`RANDOM}};
  _T_2103_re = _RAND_3830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3831 = {1{`RANDOM}};
  _T_2103_im = _RAND_3831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3832 = {1{`RANDOM}};
  _T_2104_re = _RAND_3832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3833 = {1{`RANDOM}};
  _T_2104_im = _RAND_3833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3834 = {1{`RANDOM}};
  _T_2105_re = _RAND_3834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3835 = {1{`RANDOM}};
  _T_2105_im = _RAND_3835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3836 = {1{`RANDOM}};
  _T_2106_re = _RAND_3836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3837 = {1{`RANDOM}};
  _T_2106_im = _RAND_3837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3838 = {1{`RANDOM}};
  _T_2107_re = _RAND_3838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3839 = {1{`RANDOM}};
  _T_2107_im = _RAND_3839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3840 = {1{`RANDOM}};
  _T_2108_re = _RAND_3840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3841 = {1{`RANDOM}};
  _T_2108_im = _RAND_3841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3842 = {1{`RANDOM}};
  _T_2109_re = _RAND_3842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3843 = {1{`RANDOM}};
  _T_2109_im = _RAND_3843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3844 = {1{`RANDOM}};
  _T_2110_re = _RAND_3844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3845 = {1{`RANDOM}};
  _T_2110_im = _RAND_3845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3846 = {1{`RANDOM}};
  _T_2111_re = _RAND_3846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3847 = {1{`RANDOM}};
  _T_2111_im = _RAND_3847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3848 = {1{`RANDOM}};
  _T_2112_re = _RAND_3848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3849 = {1{`RANDOM}};
  _T_2112_im = _RAND_3849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3850 = {1{`RANDOM}};
  _T_2113_re = _RAND_3850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3851 = {1{`RANDOM}};
  _T_2113_im = _RAND_3851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3852 = {1{`RANDOM}};
  _T_2114_re = _RAND_3852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3853 = {1{`RANDOM}};
  _T_2114_im = _RAND_3853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3854 = {1{`RANDOM}};
  _T_2115_re = _RAND_3854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3855 = {1{`RANDOM}};
  _T_2115_im = _RAND_3855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3856 = {1{`RANDOM}};
  _T_2116_re = _RAND_3856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3857 = {1{`RANDOM}};
  _T_2116_im = _RAND_3857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3858 = {1{`RANDOM}};
  _T_2117_re = _RAND_3858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3859 = {1{`RANDOM}};
  _T_2117_im = _RAND_3859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3860 = {1{`RANDOM}};
  _T_2118_re = _RAND_3860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3861 = {1{`RANDOM}};
  _T_2118_im = _RAND_3861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3862 = {1{`RANDOM}};
  _T_2119_re = _RAND_3862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3863 = {1{`RANDOM}};
  _T_2119_im = _RAND_3863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3864 = {1{`RANDOM}};
  _T_2120_re = _RAND_3864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3865 = {1{`RANDOM}};
  _T_2120_im = _RAND_3865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3866 = {1{`RANDOM}};
  _T_2121_re = _RAND_3866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3867 = {1{`RANDOM}};
  _T_2121_im = _RAND_3867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3868 = {1{`RANDOM}};
  _T_2122_re = _RAND_3868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3869 = {1{`RANDOM}};
  _T_2122_im = _RAND_3869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3870 = {1{`RANDOM}};
  _T_2123_re = _RAND_3870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3871 = {1{`RANDOM}};
  _T_2123_im = _RAND_3871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3872 = {1{`RANDOM}};
  _T_2124_re = _RAND_3872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3873 = {1{`RANDOM}};
  _T_2124_im = _RAND_3873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3874 = {1{`RANDOM}};
  _T_2125_re = _RAND_3874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3875 = {1{`RANDOM}};
  _T_2125_im = _RAND_3875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3876 = {1{`RANDOM}};
  _T_2126_re = _RAND_3876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3877 = {1{`RANDOM}};
  _T_2126_im = _RAND_3877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3878 = {1{`RANDOM}};
  _T_2127_re = _RAND_3878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3879 = {1{`RANDOM}};
  _T_2127_im = _RAND_3879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3880 = {1{`RANDOM}};
  _T_2128_re = _RAND_3880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3881 = {1{`RANDOM}};
  _T_2128_im = _RAND_3881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3882 = {1{`RANDOM}};
  _T_2129_re = _RAND_3882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3883 = {1{`RANDOM}};
  _T_2129_im = _RAND_3883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3884 = {1{`RANDOM}};
  _T_2130_re = _RAND_3884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3885 = {1{`RANDOM}};
  _T_2130_im = _RAND_3885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3886 = {1{`RANDOM}};
  _T_2131_re = _RAND_3886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3887 = {1{`RANDOM}};
  _T_2131_im = _RAND_3887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3888 = {1{`RANDOM}};
  _T_2132_re = _RAND_3888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3889 = {1{`RANDOM}};
  _T_2132_im = _RAND_3889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3890 = {1{`RANDOM}};
  _T_2133_re = _RAND_3890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3891 = {1{`RANDOM}};
  _T_2133_im = _RAND_3891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3892 = {1{`RANDOM}};
  _T_2134_re = _RAND_3892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3893 = {1{`RANDOM}};
  _T_2134_im = _RAND_3893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3894 = {1{`RANDOM}};
  _T_2135_re = _RAND_3894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3895 = {1{`RANDOM}};
  _T_2135_im = _RAND_3895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3896 = {1{`RANDOM}};
  _T_2136_re = _RAND_3896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3897 = {1{`RANDOM}};
  _T_2136_im = _RAND_3897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3898 = {1{`RANDOM}};
  _T_2137_re = _RAND_3898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3899 = {1{`RANDOM}};
  _T_2137_im = _RAND_3899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3900 = {1{`RANDOM}};
  _T_2138_re = _RAND_3900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3901 = {1{`RANDOM}};
  _T_2138_im = _RAND_3901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3902 = {1{`RANDOM}};
  _T_2139_re = _RAND_3902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3903 = {1{`RANDOM}};
  _T_2139_im = _RAND_3903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3904 = {1{`RANDOM}};
  _T_2140_re = _RAND_3904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3905 = {1{`RANDOM}};
  _T_2140_im = _RAND_3905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3906 = {1{`RANDOM}};
  _T_2141_re = _RAND_3906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3907 = {1{`RANDOM}};
  _T_2141_im = _RAND_3907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3908 = {1{`RANDOM}};
  _T_2142_re = _RAND_3908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3909 = {1{`RANDOM}};
  _T_2142_im = _RAND_3909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3910 = {1{`RANDOM}};
  _T_2143_re = _RAND_3910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3911 = {1{`RANDOM}};
  _T_2143_im = _RAND_3911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3912 = {1{`RANDOM}};
  _T_2144_re = _RAND_3912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3913 = {1{`RANDOM}};
  _T_2144_im = _RAND_3913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3914 = {1{`RANDOM}};
  _T_2145_re = _RAND_3914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3915 = {1{`RANDOM}};
  _T_2145_im = _RAND_3915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3916 = {1{`RANDOM}};
  _T_2146_re = _RAND_3916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3917 = {1{`RANDOM}};
  _T_2146_im = _RAND_3917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3918 = {1{`RANDOM}};
  _T_2147_re = _RAND_3918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3919 = {1{`RANDOM}};
  _T_2147_im = _RAND_3919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3920 = {1{`RANDOM}};
  _T_2148_re = _RAND_3920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3921 = {1{`RANDOM}};
  _T_2148_im = _RAND_3921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3922 = {1{`RANDOM}};
  _T_2149_re = _RAND_3922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3923 = {1{`RANDOM}};
  _T_2149_im = _RAND_3923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3924 = {1{`RANDOM}};
  _T_2150_re = _RAND_3924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3925 = {1{`RANDOM}};
  _T_2150_im = _RAND_3925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3926 = {1{`RANDOM}};
  _T_2151_re = _RAND_3926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3927 = {1{`RANDOM}};
  _T_2151_im = _RAND_3927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3928 = {1{`RANDOM}};
  _T_2152_re = _RAND_3928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3929 = {1{`RANDOM}};
  _T_2152_im = _RAND_3929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3930 = {1{`RANDOM}};
  _T_2153_re = _RAND_3930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3931 = {1{`RANDOM}};
  _T_2153_im = _RAND_3931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3932 = {1{`RANDOM}};
  _T_2154_re = _RAND_3932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3933 = {1{`RANDOM}};
  _T_2154_im = _RAND_3933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3934 = {1{`RANDOM}};
  _T_2155_re = _RAND_3934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3935 = {1{`RANDOM}};
  _T_2155_im = _RAND_3935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3936 = {1{`RANDOM}};
  _T_2156_re = _RAND_3936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3937 = {1{`RANDOM}};
  _T_2156_im = _RAND_3937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3938 = {1{`RANDOM}};
  _T_2157_re = _RAND_3938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3939 = {1{`RANDOM}};
  _T_2157_im = _RAND_3939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3940 = {1{`RANDOM}};
  _T_2158_re = _RAND_3940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3941 = {1{`RANDOM}};
  _T_2158_im = _RAND_3941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3942 = {1{`RANDOM}};
  _T_2159_re = _RAND_3942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3943 = {1{`RANDOM}};
  _T_2159_im = _RAND_3943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3944 = {1{`RANDOM}};
  _T_2160_re = _RAND_3944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3945 = {1{`RANDOM}};
  _T_2160_im = _RAND_3945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3946 = {1{`RANDOM}};
  _T_2161_re = _RAND_3946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3947 = {1{`RANDOM}};
  _T_2161_im = _RAND_3947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3948 = {1{`RANDOM}};
  _T_2162_re = _RAND_3948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3949 = {1{`RANDOM}};
  _T_2162_im = _RAND_3949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3950 = {1{`RANDOM}};
  _T_2163_re = _RAND_3950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3951 = {1{`RANDOM}};
  _T_2163_im = _RAND_3951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3952 = {1{`RANDOM}};
  _T_2164_re = _RAND_3952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3953 = {1{`RANDOM}};
  _T_2164_im = _RAND_3953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3954 = {1{`RANDOM}};
  _T_2165_re = _RAND_3954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3955 = {1{`RANDOM}};
  _T_2165_im = _RAND_3955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3956 = {1{`RANDOM}};
  _T_2166_re = _RAND_3956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3957 = {1{`RANDOM}};
  _T_2166_im = _RAND_3957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3958 = {1{`RANDOM}};
  _T_2167_re = _RAND_3958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3959 = {1{`RANDOM}};
  _T_2167_im = _RAND_3959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3960 = {1{`RANDOM}};
  _T_2168_re = _RAND_3960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3961 = {1{`RANDOM}};
  _T_2168_im = _RAND_3961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3962 = {1{`RANDOM}};
  _T_2169_re = _RAND_3962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3963 = {1{`RANDOM}};
  _T_2169_im = _RAND_3963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3964 = {1{`RANDOM}};
  _T_2170_re = _RAND_3964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3965 = {1{`RANDOM}};
  _T_2170_im = _RAND_3965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3966 = {1{`RANDOM}};
  _T_2171_re = _RAND_3966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3967 = {1{`RANDOM}};
  _T_2171_im = _RAND_3967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3968 = {1{`RANDOM}};
  _T_2172_re = _RAND_3968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3969 = {1{`RANDOM}};
  _T_2172_im = _RAND_3969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3970 = {1{`RANDOM}};
  _T_2173_re = _RAND_3970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3971 = {1{`RANDOM}};
  _T_2173_im = _RAND_3971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3972 = {1{`RANDOM}};
  _T_2174_re = _RAND_3972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3973 = {1{`RANDOM}};
  _T_2174_im = _RAND_3973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3974 = {1{`RANDOM}};
  _T_2175_re = _RAND_3974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3975 = {1{`RANDOM}};
  _T_2175_im = _RAND_3975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3976 = {1{`RANDOM}};
  _T_2176_re = _RAND_3976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3977 = {1{`RANDOM}};
  _T_2176_im = _RAND_3977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3978 = {1{`RANDOM}};
  _T_2177_re = _RAND_3978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3979 = {1{`RANDOM}};
  _T_2177_im = _RAND_3979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3980 = {1{`RANDOM}};
  _T_2178_re = _RAND_3980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3981 = {1{`RANDOM}};
  _T_2178_im = _RAND_3981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3982 = {1{`RANDOM}};
  _T_2179_re = _RAND_3982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3983 = {1{`RANDOM}};
  _T_2179_im = _RAND_3983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3984 = {1{`RANDOM}};
  _T_2180_re = _RAND_3984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3985 = {1{`RANDOM}};
  _T_2180_im = _RAND_3985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3986 = {1{`RANDOM}};
  _T_2181_re = _RAND_3986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3987 = {1{`RANDOM}};
  _T_2181_im = _RAND_3987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3988 = {1{`RANDOM}};
  _T_2182_re = _RAND_3988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3989 = {1{`RANDOM}};
  _T_2182_im = _RAND_3989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3990 = {1{`RANDOM}};
  _T_2183_re = _RAND_3990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3991 = {1{`RANDOM}};
  _T_2183_im = _RAND_3991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3992 = {1{`RANDOM}};
  _T_2184_re = _RAND_3992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3993 = {1{`RANDOM}};
  _T_2184_im = _RAND_3993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3994 = {1{`RANDOM}};
  _T_2185_re = _RAND_3994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3995 = {1{`RANDOM}};
  _T_2185_im = _RAND_3995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3996 = {1{`RANDOM}};
  _T_2186_re = _RAND_3996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3997 = {1{`RANDOM}};
  _T_2186_im = _RAND_3997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3998 = {1{`RANDOM}};
  _T_2187_re = _RAND_3998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3999 = {1{`RANDOM}};
  _T_2187_im = _RAND_3999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4000 = {1{`RANDOM}};
  _T_2188_re = _RAND_4000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4001 = {1{`RANDOM}};
  _T_2188_im = _RAND_4001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4002 = {1{`RANDOM}};
  _T_2189_re = _RAND_4002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4003 = {1{`RANDOM}};
  _T_2189_im = _RAND_4003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4004 = {1{`RANDOM}};
  _T_2190_re = _RAND_4004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4005 = {1{`RANDOM}};
  _T_2190_im = _RAND_4005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4006 = {1{`RANDOM}};
  _T_2191_re = _RAND_4006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4007 = {1{`RANDOM}};
  _T_2191_im = _RAND_4007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4008 = {1{`RANDOM}};
  _T_2192_re = _RAND_4008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4009 = {1{`RANDOM}};
  _T_2192_im = _RAND_4009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4010 = {1{`RANDOM}};
  _T_2193_re = _RAND_4010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4011 = {1{`RANDOM}};
  _T_2193_im = _RAND_4011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4012 = {1{`RANDOM}};
  _T_2194_re = _RAND_4012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4013 = {1{`RANDOM}};
  _T_2194_im = _RAND_4013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4014 = {1{`RANDOM}};
  _T_2195_re = _RAND_4014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4015 = {1{`RANDOM}};
  _T_2195_im = _RAND_4015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4016 = {1{`RANDOM}};
  _T_2196_re = _RAND_4016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4017 = {1{`RANDOM}};
  _T_2196_im = _RAND_4017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4018 = {1{`RANDOM}};
  _T_2197_re = _RAND_4018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4019 = {1{`RANDOM}};
  _T_2197_im = _RAND_4019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4020 = {1{`RANDOM}};
  _T_2198_re = _RAND_4020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4021 = {1{`RANDOM}};
  _T_2198_im = _RAND_4021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4022 = {1{`RANDOM}};
  _T_2199_re = _RAND_4022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4023 = {1{`RANDOM}};
  _T_2199_im = _RAND_4023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4024 = {1{`RANDOM}};
  _T_2200_re = _RAND_4024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4025 = {1{`RANDOM}};
  _T_2200_im = _RAND_4025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4026 = {1{`RANDOM}};
  _T_2201_re = _RAND_4026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4027 = {1{`RANDOM}};
  _T_2201_im = _RAND_4027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4028 = {1{`RANDOM}};
  _T_2202_re = _RAND_4028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4029 = {1{`RANDOM}};
  _T_2202_im = _RAND_4029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4030 = {1{`RANDOM}};
  _T_2203_re = _RAND_4030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4031 = {1{`RANDOM}};
  _T_2203_im = _RAND_4031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4032 = {1{`RANDOM}};
  _T_2204_re = _RAND_4032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4033 = {1{`RANDOM}};
  _T_2204_im = _RAND_4033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4034 = {1{`RANDOM}};
  _T_2205_re = _RAND_4034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4035 = {1{`RANDOM}};
  _T_2205_im = _RAND_4035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4036 = {1{`RANDOM}};
  _T_2206_re = _RAND_4036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4037 = {1{`RANDOM}};
  _T_2206_im = _RAND_4037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4038 = {1{`RANDOM}};
  _T_2207_re = _RAND_4038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4039 = {1{`RANDOM}};
  _T_2207_im = _RAND_4039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4040 = {1{`RANDOM}};
  _T_2208_re = _RAND_4040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4041 = {1{`RANDOM}};
  _T_2208_im = _RAND_4041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4042 = {1{`RANDOM}};
  _T_2209_re = _RAND_4042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4043 = {1{`RANDOM}};
  _T_2209_im = _RAND_4043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4044 = {1{`RANDOM}};
  _T_2210_re = _RAND_4044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4045 = {1{`RANDOM}};
  _T_2210_im = _RAND_4045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4046 = {1{`RANDOM}};
  _T_2211_re = _RAND_4046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4047 = {1{`RANDOM}};
  _T_2211_im = _RAND_4047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4048 = {1{`RANDOM}};
  _T_2212_re = _RAND_4048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4049 = {1{`RANDOM}};
  _T_2212_im = _RAND_4049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4050 = {1{`RANDOM}};
  _T_2213_re = _RAND_4050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4051 = {1{`RANDOM}};
  _T_2213_im = _RAND_4051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4052 = {1{`RANDOM}};
  _T_2214_re = _RAND_4052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4053 = {1{`RANDOM}};
  _T_2214_im = _RAND_4053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4054 = {1{`RANDOM}};
  _T_2215_re = _RAND_4054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4055 = {1{`RANDOM}};
  _T_2215_im = _RAND_4055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4056 = {1{`RANDOM}};
  _T_2216_re = _RAND_4056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4057 = {1{`RANDOM}};
  _T_2216_im = _RAND_4057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4058 = {1{`RANDOM}};
  _T_2217_re = _RAND_4058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4059 = {1{`RANDOM}};
  _T_2217_im = _RAND_4059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4060 = {1{`RANDOM}};
  _T_2218_re = _RAND_4060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4061 = {1{`RANDOM}};
  _T_2218_im = _RAND_4061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4062 = {1{`RANDOM}};
  _T_2219_re = _RAND_4062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4063 = {1{`RANDOM}};
  _T_2219_im = _RAND_4063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4064 = {1{`RANDOM}};
  _T_2220_re = _RAND_4064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4065 = {1{`RANDOM}};
  _T_2220_im = _RAND_4065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4066 = {1{`RANDOM}};
  _T_2221_re = _RAND_4066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4067 = {1{`RANDOM}};
  _T_2221_im = _RAND_4067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4068 = {1{`RANDOM}};
  _T_2222_re = _RAND_4068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4069 = {1{`RANDOM}};
  _T_2222_im = _RAND_4069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4070 = {1{`RANDOM}};
  _T_2223_re = _RAND_4070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4071 = {1{`RANDOM}};
  _T_2223_im = _RAND_4071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4072 = {1{`RANDOM}};
  _T_2224_re = _RAND_4072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4073 = {1{`RANDOM}};
  _T_2224_im = _RAND_4073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4074 = {1{`RANDOM}};
  _T_2225_re = _RAND_4074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4075 = {1{`RANDOM}};
  _T_2225_im = _RAND_4075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4076 = {1{`RANDOM}};
  _T_2226_re = _RAND_4076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4077 = {1{`RANDOM}};
  _T_2226_im = _RAND_4077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4078 = {1{`RANDOM}};
  _T_2227_re = _RAND_4078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4079 = {1{`RANDOM}};
  _T_2227_im = _RAND_4079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4080 = {1{`RANDOM}};
  _T_2228_re = _RAND_4080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4081 = {1{`RANDOM}};
  _T_2228_im = _RAND_4081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4082 = {1{`RANDOM}};
  _T_2229_re = _RAND_4082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4083 = {1{`RANDOM}};
  _T_2229_im = _RAND_4083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4084 = {1{`RANDOM}};
  _T_2230_re = _RAND_4084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4085 = {1{`RANDOM}};
  _T_2230_im = _RAND_4085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4086 = {1{`RANDOM}};
  _T_2231_re = _RAND_4086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4087 = {1{`RANDOM}};
  _T_2231_im = _RAND_4087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4088 = {1{`RANDOM}};
  _T_2232_re = _RAND_4088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4089 = {1{`RANDOM}};
  _T_2232_im = _RAND_4089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4090 = {1{`RANDOM}};
  _T_2233_re = _RAND_4090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4091 = {1{`RANDOM}};
  _T_2233_im = _RAND_4091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4092 = {1{`RANDOM}};
  _T_2234_re = _RAND_4092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4093 = {1{`RANDOM}};
  _T_2234_im = _RAND_4093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4094 = {1{`RANDOM}};
  _T_2235_re = _RAND_4094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4095 = {1{`RANDOM}};
  _T_2235_im = _RAND_4095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4096 = {1{`RANDOM}};
  _T_2236_re = _RAND_4096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4097 = {1{`RANDOM}};
  _T_2236_im = _RAND_4097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4098 = {1{`RANDOM}};
  _T_2239_re = _RAND_4098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4099 = {1{`RANDOM}};
  _T_2239_im = _RAND_4099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4100 = {1{`RANDOM}};
  _T_2240_re = _RAND_4100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4101 = {1{`RANDOM}};
  _T_2240_im = _RAND_4101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4102 = {1{`RANDOM}};
  _T_2241_re = _RAND_4102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4103 = {1{`RANDOM}};
  _T_2241_im = _RAND_4103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4104 = {1{`RANDOM}};
  _T_2242_re = _RAND_4104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4105 = {1{`RANDOM}};
  _T_2242_im = _RAND_4105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4106 = {1{`RANDOM}};
  _T_2243_re = _RAND_4106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4107 = {1{`RANDOM}};
  _T_2243_im = _RAND_4107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4108 = {1{`RANDOM}};
  _T_2244_re = _RAND_4108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4109 = {1{`RANDOM}};
  _T_2244_im = _RAND_4109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4110 = {1{`RANDOM}};
  _T_2245_re = _RAND_4110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4111 = {1{`RANDOM}};
  _T_2245_im = _RAND_4111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4112 = {1{`RANDOM}};
  _T_2246_re = _RAND_4112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4113 = {1{`RANDOM}};
  _T_2246_im = _RAND_4113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4114 = {1{`RANDOM}};
  _T_2247_re = _RAND_4114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4115 = {1{`RANDOM}};
  _T_2247_im = _RAND_4115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4116 = {1{`RANDOM}};
  _T_2248_re = _RAND_4116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4117 = {1{`RANDOM}};
  _T_2248_im = _RAND_4117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4118 = {1{`RANDOM}};
  _T_2249_re = _RAND_4118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4119 = {1{`RANDOM}};
  _T_2249_im = _RAND_4119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4120 = {1{`RANDOM}};
  _T_2250_re = _RAND_4120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4121 = {1{`RANDOM}};
  _T_2250_im = _RAND_4121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4122 = {1{`RANDOM}};
  _T_2251_re = _RAND_4122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4123 = {1{`RANDOM}};
  _T_2251_im = _RAND_4123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4124 = {1{`RANDOM}};
  _T_2252_re = _RAND_4124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4125 = {1{`RANDOM}};
  _T_2252_im = _RAND_4125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4126 = {1{`RANDOM}};
  _T_2253_re = _RAND_4126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4127 = {1{`RANDOM}};
  _T_2253_im = _RAND_4127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4128 = {1{`RANDOM}};
  _T_2254_re = _RAND_4128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4129 = {1{`RANDOM}};
  _T_2254_im = _RAND_4129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4130 = {1{`RANDOM}};
  _T_2255_re = _RAND_4130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4131 = {1{`RANDOM}};
  _T_2255_im = _RAND_4131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4132 = {1{`RANDOM}};
  _T_2256_re = _RAND_4132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4133 = {1{`RANDOM}};
  _T_2256_im = _RAND_4133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4134 = {1{`RANDOM}};
  _T_2257_re = _RAND_4134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4135 = {1{`RANDOM}};
  _T_2257_im = _RAND_4135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4136 = {1{`RANDOM}};
  _T_2258_re = _RAND_4136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4137 = {1{`RANDOM}};
  _T_2258_im = _RAND_4137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4138 = {1{`RANDOM}};
  _T_2259_re = _RAND_4138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4139 = {1{`RANDOM}};
  _T_2259_im = _RAND_4139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4140 = {1{`RANDOM}};
  _T_2260_re = _RAND_4140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4141 = {1{`RANDOM}};
  _T_2260_im = _RAND_4141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4142 = {1{`RANDOM}};
  _T_2261_re = _RAND_4142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4143 = {1{`RANDOM}};
  _T_2261_im = _RAND_4143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4144 = {1{`RANDOM}};
  _T_2262_re = _RAND_4144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4145 = {1{`RANDOM}};
  _T_2262_im = _RAND_4145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4146 = {1{`RANDOM}};
  _T_2263_re = _RAND_4146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4147 = {1{`RANDOM}};
  _T_2263_im = _RAND_4147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4148 = {1{`RANDOM}};
  _T_2264_re = _RAND_4148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4149 = {1{`RANDOM}};
  _T_2264_im = _RAND_4149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4150 = {1{`RANDOM}};
  _T_2265_re = _RAND_4150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4151 = {1{`RANDOM}};
  _T_2265_im = _RAND_4151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4152 = {1{`RANDOM}};
  _T_2266_re = _RAND_4152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4153 = {1{`RANDOM}};
  _T_2266_im = _RAND_4153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4154 = {1{`RANDOM}};
  _T_2267_re = _RAND_4154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4155 = {1{`RANDOM}};
  _T_2267_im = _RAND_4155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4156 = {1{`RANDOM}};
  _T_2268_re = _RAND_4156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4157 = {1{`RANDOM}};
  _T_2268_im = _RAND_4157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4158 = {1{`RANDOM}};
  _T_2269_re = _RAND_4158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4159 = {1{`RANDOM}};
  _T_2269_im = _RAND_4159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4160 = {1{`RANDOM}};
  _T_2270_re = _RAND_4160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4161 = {1{`RANDOM}};
  _T_2270_im = _RAND_4161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4162 = {1{`RANDOM}};
  _T_2271_re = _RAND_4162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4163 = {1{`RANDOM}};
  _T_2271_im = _RAND_4163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4164 = {1{`RANDOM}};
  _T_2272_re = _RAND_4164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4165 = {1{`RANDOM}};
  _T_2272_im = _RAND_4165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4166 = {1{`RANDOM}};
  _T_2273_re = _RAND_4166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4167 = {1{`RANDOM}};
  _T_2273_im = _RAND_4167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4168 = {1{`RANDOM}};
  _T_2274_re = _RAND_4168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4169 = {1{`RANDOM}};
  _T_2274_im = _RAND_4169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4170 = {1{`RANDOM}};
  _T_2275_re = _RAND_4170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4171 = {1{`RANDOM}};
  _T_2275_im = _RAND_4171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4172 = {1{`RANDOM}};
  _T_2276_re = _RAND_4172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4173 = {1{`RANDOM}};
  _T_2276_im = _RAND_4173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4174 = {1{`RANDOM}};
  _T_2277_re = _RAND_4174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4175 = {1{`RANDOM}};
  _T_2277_im = _RAND_4175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4176 = {1{`RANDOM}};
  _T_2278_re = _RAND_4176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4177 = {1{`RANDOM}};
  _T_2278_im = _RAND_4177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4178 = {1{`RANDOM}};
  _T_2279_re = _RAND_4178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4179 = {1{`RANDOM}};
  _T_2279_im = _RAND_4179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4180 = {1{`RANDOM}};
  _T_2280_re = _RAND_4180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4181 = {1{`RANDOM}};
  _T_2280_im = _RAND_4181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4182 = {1{`RANDOM}};
  _T_2281_re = _RAND_4182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4183 = {1{`RANDOM}};
  _T_2281_im = _RAND_4183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4184 = {1{`RANDOM}};
  _T_2282_re = _RAND_4184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4185 = {1{`RANDOM}};
  _T_2282_im = _RAND_4185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4186 = {1{`RANDOM}};
  _T_2283_re = _RAND_4186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4187 = {1{`RANDOM}};
  _T_2283_im = _RAND_4187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4188 = {1{`RANDOM}};
  _T_2284_re = _RAND_4188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4189 = {1{`RANDOM}};
  _T_2284_im = _RAND_4189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4190 = {1{`RANDOM}};
  _T_2285_re = _RAND_4190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4191 = {1{`RANDOM}};
  _T_2285_im = _RAND_4191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4192 = {1{`RANDOM}};
  _T_2286_re = _RAND_4192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4193 = {1{`RANDOM}};
  _T_2286_im = _RAND_4193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4194 = {1{`RANDOM}};
  _T_2287_re = _RAND_4194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4195 = {1{`RANDOM}};
  _T_2287_im = _RAND_4195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4196 = {1{`RANDOM}};
  _T_2288_re = _RAND_4196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4197 = {1{`RANDOM}};
  _T_2288_im = _RAND_4197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4198 = {1{`RANDOM}};
  _T_2289_re = _RAND_4198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4199 = {1{`RANDOM}};
  _T_2289_im = _RAND_4199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4200 = {1{`RANDOM}};
  _T_2290_re = _RAND_4200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4201 = {1{`RANDOM}};
  _T_2290_im = _RAND_4201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4202 = {1{`RANDOM}};
  _T_2291_re = _RAND_4202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4203 = {1{`RANDOM}};
  _T_2291_im = _RAND_4203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4204 = {1{`RANDOM}};
  _T_2292_re = _RAND_4204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4205 = {1{`RANDOM}};
  _T_2292_im = _RAND_4205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4206 = {1{`RANDOM}};
  _T_2293_re = _RAND_4206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4207 = {1{`RANDOM}};
  _T_2293_im = _RAND_4207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4208 = {1{`RANDOM}};
  _T_2294_re = _RAND_4208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4209 = {1{`RANDOM}};
  _T_2294_im = _RAND_4209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4210 = {1{`RANDOM}};
  _T_2295_re = _RAND_4210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4211 = {1{`RANDOM}};
  _T_2295_im = _RAND_4211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4212 = {1{`RANDOM}};
  _T_2296_re = _RAND_4212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4213 = {1{`RANDOM}};
  _T_2296_im = _RAND_4213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4214 = {1{`RANDOM}};
  _T_2297_re = _RAND_4214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4215 = {1{`RANDOM}};
  _T_2297_im = _RAND_4215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4216 = {1{`RANDOM}};
  _T_2298_re = _RAND_4216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4217 = {1{`RANDOM}};
  _T_2298_im = _RAND_4217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4218 = {1{`RANDOM}};
  _T_2299_re = _RAND_4218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4219 = {1{`RANDOM}};
  _T_2299_im = _RAND_4219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4220 = {1{`RANDOM}};
  _T_2300_re = _RAND_4220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4221 = {1{`RANDOM}};
  _T_2300_im = _RAND_4221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4222 = {1{`RANDOM}};
  _T_2301_re = _RAND_4222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4223 = {1{`RANDOM}};
  _T_2301_im = _RAND_4223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4224 = {1{`RANDOM}};
  _T_2302_re = _RAND_4224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4225 = {1{`RANDOM}};
  _T_2302_im = _RAND_4225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4226 = {1{`RANDOM}};
  _T_2303_re = _RAND_4226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4227 = {1{`RANDOM}};
  _T_2303_im = _RAND_4227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4228 = {1{`RANDOM}};
  _T_2304_re = _RAND_4228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4229 = {1{`RANDOM}};
  _T_2304_im = _RAND_4229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4230 = {1{`RANDOM}};
  _T_2305_re = _RAND_4230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4231 = {1{`RANDOM}};
  _T_2305_im = _RAND_4231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4232 = {1{`RANDOM}};
  _T_2306_re = _RAND_4232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4233 = {1{`RANDOM}};
  _T_2306_im = _RAND_4233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4234 = {1{`RANDOM}};
  _T_2307_re = _RAND_4234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4235 = {1{`RANDOM}};
  _T_2307_im = _RAND_4235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4236 = {1{`RANDOM}};
  _T_2308_re = _RAND_4236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4237 = {1{`RANDOM}};
  _T_2308_im = _RAND_4237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4238 = {1{`RANDOM}};
  _T_2309_re = _RAND_4238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4239 = {1{`RANDOM}};
  _T_2309_im = _RAND_4239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4240 = {1{`RANDOM}};
  _T_2310_re = _RAND_4240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4241 = {1{`RANDOM}};
  _T_2310_im = _RAND_4241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4242 = {1{`RANDOM}};
  _T_2311_re = _RAND_4242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4243 = {1{`RANDOM}};
  _T_2311_im = _RAND_4243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4244 = {1{`RANDOM}};
  _T_2312_re = _RAND_4244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4245 = {1{`RANDOM}};
  _T_2312_im = _RAND_4245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4246 = {1{`RANDOM}};
  _T_2313_re = _RAND_4246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4247 = {1{`RANDOM}};
  _T_2313_im = _RAND_4247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4248 = {1{`RANDOM}};
  _T_2314_re = _RAND_4248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4249 = {1{`RANDOM}};
  _T_2314_im = _RAND_4249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4250 = {1{`RANDOM}};
  _T_2315_re = _RAND_4250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4251 = {1{`RANDOM}};
  _T_2315_im = _RAND_4251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4252 = {1{`RANDOM}};
  _T_2316_re = _RAND_4252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4253 = {1{`RANDOM}};
  _T_2316_im = _RAND_4253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4254 = {1{`RANDOM}};
  _T_2317_re = _RAND_4254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4255 = {1{`RANDOM}};
  _T_2317_im = _RAND_4255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4256 = {1{`RANDOM}};
  _T_2318_re = _RAND_4256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4257 = {1{`RANDOM}};
  _T_2318_im = _RAND_4257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4258 = {1{`RANDOM}};
  _T_2319_re = _RAND_4258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4259 = {1{`RANDOM}};
  _T_2319_im = _RAND_4259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4260 = {1{`RANDOM}};
  _T_2320_re = _RAND_4260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4261 = {1{`RANDOM}};
  _T_2320_im = _RAND_4261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4262 = {1{`RANDOM}};
  _T_2321_re = _RAND_4262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4263 = {1{`RANDOM}};
  _T_2321_im = _RAND_4263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4264 = {1{`RANDOM}};
  _T_2322_re = _RAND_4264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4265 = {1{`RANDOM}};
  _T_2322_im = _RAND_4265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4266 = {1{`RANDOM}};
  _T_2323_re = _RAND_4266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4267 = {1{`RANDOM}};
  _T_2323_im = _RAND_4267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4268 = {1{`RANDOM}};
  _T_2324_re = _RAND_4268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4269 = {1{`RANDOM}};
  _T_2324_im = _RAND_4269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4270 = {1{`RANDOM}};
  _T_2325_re = _RAND_4270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4271 = {1{`RANDOM}};
  _T_2325_im = _RAND_4271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4272 = {1{`RANDOM}};
  _T_2326_re = _RAND_4272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4273 = {1{`RANDOM}};
  _T_2326_im = _RAND_4273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4274 = {1{`RANDOM}};
  _T_2327_re = _RAND_4274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4275 = {1{`RANDOM}};
  _T_2327_im = _RAND_4275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4276 = {1{`RANDOM}};
  _T_2328_re = _RAND_4276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4277 = {1{`RANDOM}};
  _T_2328_im = _RAND_4277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4278 = {1{`RANDOM}};
  _T_2329_re = _RAND_4278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4279 = {1{`RANDOM}};
  _T_2329_im = _RAND_4279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4280 = {1{`RANDOM}};
  _T_2330_re = _RAND_4280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4281 = {1{`RANDOM}};
  _T_2330_im = _RAND_4281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4282 = {1{`RANDOM}};
  _T_2331_re = _RAND_4282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4283 = {1{`RANDOM}};
  _T_2331_im = _RAND_4283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4284 = {1{`RANDOM}};
  _T_2332_re = _RAND_4284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4285 = {1{`RANDOM}};
  _T_2332_im = _RAND_4285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4286 = {1{`RANDOM}};
  _T_2333_re = _RAND_4286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4287 = {1{`RANDOM}};
  _T_2333_im = _RAND_4287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4288 = {1{`RANDOM}};
  _T_2334_re = _RAND_4288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4289 = {1{`RANDOM}};
  _T_2334_im = _RAND_4289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4290 = {1{`RANDOM}};
  _T_2335_re = _RAND_4290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4291 = {1{`RANDOM}};
  _T_2335_im = _RAND_4291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4292 = {1{`RANDOM}};
  _T_2336_re = _RAND_4292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4293 = {1{`RANDOM}};
  _T_2336_im = _RAND_4293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4294 = {1{`RANDOM}};
  _T_2337_re = _RAND_4294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4295 = {1{`RANDOM}};
  _T_2337_im = _RAND_4295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4296 = {1{`RANDOM}};
  _T_2338_re = _RAND_4296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4297 = {1{`RANDOM}};
  _T_2338_im = _RAND_4297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4298 = {1{`RANDOM}};
  _T_2339_re = _RAND_4298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4299 = {1{`RANDOM}};
  _T_2339_im = _RAND_4299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4300 = {1{`RANDOM}};
  _T_2340_re = _RAND_4300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4301 = {1{`RANDOM}};
  _T_2340_im = _RAND_4301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4302 = {1{`RANDOM}};
  _T_2341_re = _RAND_4302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4303 = {1{`RANDOM}};
  _T_2341_im = _RAND_4303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4304 = {1{`RANDOM}};
  _T_2342_re = _RAND_4304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4305 = {1{`RANDOM}};
  _T_2342_im = _RAND_4305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4306 = {1{`RANDOM}};
  _T_2343_re = _RAND_4306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4307 = {1{`RANDOM}};
  _T_2343_im = _RAND_4307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4308 = {1{`RANDOM}};
  _T_2344_re = _RAND_4308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4309 = {1{`RANDOM}};
  _T_2344_im = _RAND_4309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4310 = {1{`RANDOM}};
  _T_2345_re = _RAND_4310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4311 = {1{`RANDOM}};
  _T_2345_im = _RAND_4311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4312 = {1{`RANDOM}};
  _T_2346_re = _RAND_4312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4313 = {1{`RANDOM}};
  _T_2346_im = _RAND_4313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4314 = {1{`RANDOM}};
  _T_2347_re = _RAND_4314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4315 = {1{`RANDOM}};
  _T_2347_im = _RAND_4315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4316 = {1{`RANDOM}};
  _T_2348_re = _RAND_4316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4317 = {1{`RANDOM}};
  _T_2348_im = _RAND_4317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4318 = {1{`RANDOM}};
  _T_2349_re = _RAND_4318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4319 = {1{`RANDOM}};
  _T_2349_im = _RAND_4319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4320 = {1{`RANDOM}};
  _T_2350_re = _RAND_4320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4321 = {1{`RANDOM}};
  _T_2350_im = _RAND_4321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4322 = {1{`RANDOM}};
  _T_2351_re = _RAND_4322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4323 = {1{`RANDOM}};
  _T_2351_im = _RAND_4323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4324 = {1{`RANDOM}};
  _T_2352_re = _RAND_4324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4325 = {1{`RANDOM}};
  _T_2352_im = _RAND_4325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4326 = {1{`RANDOM}};
  _T_2353_re = _RAND_4326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4327 = {1{`RANDOM}};
  _T_2353_im = _RAND_4327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4328 = {1{`RANDOM}};
  _T_2354_re = _RAND_4328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4329 = {1{`RANDOM}};
  _T_2354_im = _RAND_4329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4330 = {1{`RANDOM}};
  _T_2355_re = _RAND_4330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4331 = {1{`RANDOM}};
  _T_2355_im = _RAND_4331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4332 = {1{`RANDOM}};
  _T_2356_re = _RAND_4332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4333 = {1{`RANDOM}};
  _T_2356_im = _RAND_4333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4334 = {1{`RANDOM}};
  _T_2357_re = _RAND_4334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4335 = {1{`RANDOM}};
  _T_2357_im = _RAND_4335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4336 = {1{`RANDOM}};
  _T_2358_re = _RAND_4336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4337 = {1{`RANDOM}};
  _T_2358_im = _RAND_4337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4338 = {1{`RANDOM}};
  _T_2359_re = _RAND_4338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4339 = {1{`RANDOM}};
  _T_2359_im = _RAND_4339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4340 = {1{`RANDOM}};
  _T_2360_re = _RAND_4340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4341 = {1{`RANDOM}};
  _T_2360_im = _RAND_4341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4342 = {1{`RANDOM}};
  _T_2361_re = _RAND_4342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4343 = {1{`RANDOM}};
  _T_2361_im = _RAND_4343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4344 = {1{`RANDOM}};
  _T_2362_re = _RAND_4344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4345 = {1{`RANDOM}};
  _T_2362_im = _RAND_4345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4346 = {1{`RANDOM}};
  _T_2363_re = _RAND_4346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4347 = {1{`RANDOM}};
  _T_2363_im = _RAND_4347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4348 = {1{`RANDOM}};
  _T_2364_re = _RAND_4348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4349 = {1{`RANDOM}};
  _T_2364_im = _RAND_4349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4350 = {1{`RANDOM}};
  _T_2365_re = _RAND_4350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4351 = {1{`RANDOM}};
  _T_2365_im = _RAND_4351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4352 = {1{`RANDOM}};
  _T_2366_re = _RAND_4352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4353 = {1{`RANDOM}};
  _T_2366_im = _RAND_4353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4354 = {1{`RANDOM}};
  _T_2367_re = _RAND_4354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4355 = {1{`RANDOM}};
  _T_2367_im = _RAND_4355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4356 = {1{`RANDOM}};
  _T_2368_re = _RAND_4356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4357 = {1{`RANDOM}};
  _T_2368_im = _RAND_4357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4358 = {1{`RANDOM}};
  _T_2369_re = _RAND_4358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4359 = {1{`RANDOM}};
  _T_2369_im = _RAND_4359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4360 = {1{`RANDOM}};
  _T_2370_re = _RAND_4360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4361 = {1{`RANDOM}};
  _T_2370_im = _RAND_4361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4362 = {1{`RANDOM}};
  _T_2371_re = _RAND_4362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4363 = {1{`RANDOM}};
  _T_2371_im = _RAND_4363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4364 = {1{`RANDOM}};
  _T_2372_re = _RAND_4364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4365 = {1{`RANDOM}};
  _T_2372_im = _RAND_4365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4366 = {1{`RANDOM}};
  _T_2373_re = _RAND_4366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4367 = {1{`RANDOM}};
  _T_2373_im = _RAND_4367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4368 = {1{`RANDOM}};
  _T_2374_re = _RAND_4368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4369 = {1{`RANDOM}};
  _T_2374_im = _RAND_4369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4370 = {1{`RANDOM}};
  _T_2375_re = _RAND_4370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4371 = {1{`RANDOM}};
  _T_2375_im = _RAND_4371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4372 = {1{`RANDOM}};
  _T_2376_re = _RAND_4372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4373 = {1{`RANDOM}};
  _T_2376_im = _RAND_4373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4374 = {1{`RANDOM}};
  _T_2377_re = _RAND_4374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4375 = {1{`RANDOM}};
  _T_2377_im = _RAND_4375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4376 = {1{`RANDOM}};
  _T_2378_re = _RAND_4376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4377 = {1{`RANDOM}};
  _T_2378_im = _RAND_4377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4378 = {1{`RANDOM}};
  _T_2379_re = _RAND_4378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4379 = {1{`RANDOM}};
  _T_2379_im = _RAND_4379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4380 = {1{`RANDOM}};
  _T_2380_re = _RAND_4380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4381 = {1{`RANDOM}};
  _T_2380_im = _RAND_4381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4382 = {1{`RANDOM}};
  _T_2381_re = _RAND_4382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4383 = {1{`RANDOM}};
  _T_2381_im = _RAND_4383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4384 = {1{`RANDOM}};
  _T_2382_re = _RAND_4384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4385 = {1{`RANDOM}};
  _T_2382_im = _RAND_4385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4386 = {1{`RANDOM}};
  _T_2383_re = _RAND_4386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4387 = {1{`RANDOM}};
  _T_2383_im = _RAND_4387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4388 = {1{`RANDOM}};
  _T_2384_re = _RAND_4388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4389 = {1{`RANDOM}};
  _T_2384_im = _RAND_4389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4390 = {1{`RANDOM}};
  _T_2385_re = _RAND_4390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4391 = {1{`RANDOM}};
  _T_2385_im = _RAND_4391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4392 = {1{`RANDOM}};
  _T_2386_re = _RAND_4392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4393 = {1{`RANDOM}};
  _T_2386_im = _RAND_4393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4394 = {1{`RANDOM}};
  _T_2387_re = _RAND_4394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4395 = {1{`RANDOM}};
  _T_2387_im = _RAND_4395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4396 = {1{`RANDOM}};
  _T_2388_re = _RAND_4396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4397 = {1{`RANDOM}};
  _T_2388_im = _RAND_4397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4398 = {1{`RANDOM}};
  _T_2389_re = _RAND_4398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4399 = {1{`RANDOM}};
  _T_2389_im = _RAND_4399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4400 = {1{`RANDOM}};
  _T_2390_re = _RAND_4400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4401 = {1{`RANDOM}};
  _T_2390_im = _RAND_4401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4402 = {1{`RANDOM}};
  _T_2391_re = _RAND_4402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4403 = {1{`RANDOM}};
  _T_2391_im = _RAND_4403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4404 = {1{`RANDOM}};
  _T_2392_re = _RAND_4404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4405 = {1{`RANDOM}};
  _T_2392_im = _RAND_4405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4406 = {1{`RANDOM}};
  _T_2393_re = _RAND_4406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4407 = {1{`RANDOM}};
  _T_2393_im = _RAND_4407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4408 = {1{`RANDOM}};
  _T_2394_re = _RAND_4408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4409 = {1{`RANDOM}};
  _T_2394_im = _RAND_4409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4410 = {1{`RANDOM}};
  _T_2395_re = _RAND_4410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4411 = {1{`RANDOM}};
  _T_2395_im = _RAND_4411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4412 = {1{`RANDOM}};
  _T_2396_re = _RAND_4412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4413 = {1{`RANDOM}};
  _T_2396_im = _RAND_4413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4414 = {1{`RANDOM}};
  _T_2397_re = _RAND_4414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4415 = {1{`RANDOM}};
  _T_2397_im = _RAND_4415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4416 = {1{`RANDOM}};
  _T_2398_re = _RAND_4416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4417 = {1{`RANDOM}};
  _T_2398_im = _RAND_4417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4418 = {1{`RANDOM}};
  _T_2399_re = _RAND_4418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4419 = {1{`RANDOM}};
  _T_2399_im = _RAND_4419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4420 = {1{`RANDOM}};
  _T_2400_re = _RAND_4420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4421 = {1{`RANDOM}};
  _T_2400_im = _RAND_4421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4422 = {1{`RANDOM}};
  _T_2401_re = _RAND_4422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4423 = {1{`RANDOM}};
  _T_2401_im = _RAND_4423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4424 = {1{`RANDOM}};
  _T_2402_re = _RAND_4424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4425 = {1{`RANDOM}};
  _T_2402_im = _RAND_4425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4426 = {1{`RANDOM}};
  _T_2403_re = _RAND_4426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4427 = {1{`RANDOM}};
  _T_2403_im = _RAND_4427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4428 = {1{`RANDOM}};
  _T_2404_re = _RAND_4428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4429 = {1{`RANDOM}};
  _T_2404_im = _RAND_4429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4430 = {1{`RANDOM}};
  _T_2405_re = _RAND_4430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4431 = {1{`RANDOM}};
  _T_2405_im = _RAND_4431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4432 = {1{`RANDOM}};
  _T_2406_re = _RAND_4432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4433 = {1{`RANDOM}};
  _T_2406_im = _RAND_4433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4434 = {1{`RANDOM}};
  _T_2407_re = _RAND_4434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4435 = {1{`RANDOM}};
  _T_2407_im = _RAND_4435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4436 = {1{`RANDOM}};
  _T_2408_re = _RAND_4436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4437 = {1{`RANDOM}};
  _T_2408_im = _RAND_4437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4438 = {1{`RANDOM}};
  _T_2409_re = _RAND_4438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4439 = {1{`RANDOM}};
  _T_2409_im = _RAND_4439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4440 = {1{`RANDOM}};
  _T_2410_re = _RAND_4440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4441 = {1{`RANDOM}};
  _T_2410_im = _RAND_4441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4442 = {1{`RANDOM}};
  _T_2411_re = _RAND_4442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4443 = {1{`RANDOM}};
  _T_2411_im = _RAND_4443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4444 = {1{`RANDOM}};
  _T_2412_re = _RAND_4444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4445 = {1{`RANDOM}};
  _T_2412_im = _RAND_4445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4446 = {1{`RANDOM}};
  _T_2413_re = _RAND_4446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4447 = {1{`RANDOM}};
  _T_2413_im = _RAND_4447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4448 = {1{`RANDOM}};
  _T_2414_re = _RAND_4448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4449 = {1{`RANDOM}};
  _T_2414_im = _RAND_4449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4450 = {1{`RANDOM}};
  _T_2415_re = _RAND_4450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4451 = {1{`RANDOM}};
  _T_2415_im = _RAND_4451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4452 = {1{`RANDOM}};
  _T_2416_re = _RAND_4452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4453 = {1{`RANDOM}};
  _T_2416_im = _RAND_4453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4454 = {1{`RANDOM}};
  _T_2417_re = _RAND_4454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4455 = {1{`RANDOM}};
  _T_2417_im = _RAND_4455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4456 = {1{`RANDOM}};
  _T_2418_re = _RAND_4456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4457 = {1{`RANDOM}};
  _T_2418_im = _RAND_4457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4458 = {1{`RANDOM}};
  _T_2419_re = _RAND_4458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4459 = {1{`RANDOM}};
  _T_2419_im = _RAND_4459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4460 = {1{`RANDOM}};
  _T_2420_re = _RAND_4460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4461 = {1{`RANDOM}};
  _T_2420_im = _RAND_4461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4462 = {1{`RANDOM}};
  _T_2421_re = _RAND_4462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4463 = {1{`RANDOM}};
  _T_2421_im = _RAND_4463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4464 = {1{`RANDOM}};
  _T_2422_re = _RAND_4464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4465 = {1{`RANDOM}};
  _T_2422_im = _RAND_4465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4466 = {1{`RANDOM}};
  _T_2423_re = _RAND_4466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4467 = {1{`RANDOM}};
  _T_2423_im = _RAND_4467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4468 = {1{`RANDOM}};
  _T_2424_re = _RAND_4468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4469 = {1{`RANDOM}};
  _T_2424_im = _RAND_4469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4470 = {1{`RANDOM}};
  _T_2425_re = _RAND_4470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4471 = {1{`RANDOM}};
  _T_2425_im = _RAND_4471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4472 = {1{`RANDOM}};
  _T_2426_re = _RAND_4472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4473 = {1{`RANDOM}};
  _T_2426_im = _RAND_4473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4474 = {1{`RANDOM}};
  _T_2427_re = _RAND_4474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4475 = {1{`RANDOM}};
  _T_2427_im = _RAND_4475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4476 = {1{`RANDOM}};
  _T_2428_re = _RAND_4476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4477 = {1{`RANDOM}};
  _T_2428_im = _RAND_4477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4478 = {1{`RANDOM}};
  _T_2429_re = _RAND_4478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4479 = {1{`RANDOM}};
  _T_2429_im = _RAND_4479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4480 = {1{`RANDOM}};
  _T_2430_re = _RAND_4480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4481 = {1{`RANDOM}};
  _T_2430_im = _RAND_4481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4482 = {1{`RANDOM}};
  _T_2431_re = _RAND_4482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4483 = {1{`RANDOM}};
  _T_2431_im = _RAND_4483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4484 = {1{`RANDOM}};
  _T_2432_re = _RAND_4484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4485 = {1{`RANDOM}};
  _T_2432_im = _RAND_4485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4486 = {1{`RANDOM}};
  _T_2433_re = _RAND_4486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4487 = {1{`RANDOM}};
  _T_2433_im = _RAND_4487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4488 = {1{`RANDOM}};
  _T_2434_re = _RAND_4488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4489 = {1{`RANDOM}};
  _T_2434_im = _RAND_4489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4490 = {1{`RANDOM}};
  _T_2435_re = _RAND_4490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4491 = {1{`RANDOM}};
  _T_2435_im = _RAND_4491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4492 = {1{`RANDOM}};
  _T_2436_re = _RAND_4492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4493 = {1{`RANDOM}};
  _T_2436_im = _RAND_4493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4494 = {1{`RANDOM}};
  _T_2437_re = _RAND_4494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4495 = {1{`RANDOM}};
  _T_2437_im = _RAND_4495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4496 = {1{`RANDOM}};
  _T_2438_re = _RAND_4496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4497 = {1{`RANDOM}};
  _T_2438_im = _RAND_4497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4498 = {1{`RANDOM}};
  _T_2439_re = _RAND_4498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4499 = {1{`RANDOM}};
  _T_2439_im = _RAND_4499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4500 = {1{`RANDOM}};
  _T_2440_re = _RAND_4500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4501 = {1{`RANDOM}};
  _T_2440_im = _RAND_4501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4502 = {1{`RANDOM}};
  _T_2441_re = _RAND_4502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4503 = {1{`RANDOM}};
  _T_2441_im = _RAND_4503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4504 = {1{`RANDOM}};
  _T_2442_re = _RAND_4504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4505 = {1{`RANDOM}};
  _T_2442_im = _RAND_4505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4506 = {1{`RANDOM}};
  _T_2443_re = _RAND_4506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4507 = {1{`RANDOM}};
  _T_2443_im = _RAND_4507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4508 = {1{`RANDOM}};
  _T_2444_re = _RAND_4508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4509 = {1{`RANDOM}};
  _T_2444_im = _RAND_4509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4510 = {1{`RANDOM}};
  _T_2445_re = _RAND_4510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4511 = {1{`RANDOM}};
  _T_2445_im = _RAND_4511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4512 = {1{`RANDOM}};
  _T_2446_re = _RAND_4512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4513 = {1{`RANDOM}};
  _T_2446_im = _RAND_4513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4514 = {1{`RANDOM}};
  _T_2447_re = _RAND_4514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4515 = {1{`RANDOM}};
  _T_2447_im = _RAND_4515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4516 = {1{`RANDOM}};
  _T_2448_re = _RAND_4516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4517 = {1{`RANDOM}};
  _T_2448_im = _RAND_4517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4518 = {1{`RANDOM}};
  _T_2449_re = _RAND_4518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4519 = {1{`RANDOM}};
  _T_2449_im = _RAND_4519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4520 = {1{`RANDOM}};
  _T_2450_re = _RAND_4520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4521 = {1{`RANDOM}};
  _T_2450_im = _RAND_4521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4522 = {1{`RANDOM}};
  _T_2451_re = _RAND_4522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4523 = {1{`RANDOM}};
  _T_2451_im = _RAND_4523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4524 = {1{`RANDOM}};
  _T_2452_re = _RAND_4524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4525 = {1{`RANDOM}};
  _T_2452_im = _RAND_4525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4526 = {1{`RANDOM}};
  _T_2453_re = _RAND_4526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4527 = {1{`RANDOM}};
  _T_2453_im = _RAND_4527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4528 = {1{`RANDOM}};
  _T_2454_re = _RAND_4528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4529 = {1{`RANDOM}};
  _T_2454_im = _RAND_4529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4530 = {1{`RANDOM}};
  _T_2455_re = _RAND_4530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4531 = {1{`RANDOM}};
  _T_2455_im = _RAND_4531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4532 = {1{`RANDOM}};
  _T_2456_re = _RAND_4532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4533 = {1{`RANDOM}};
  _T_2456_im = _RAND_4533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4534 = {1{`RANDOM}};
  _T_2457_re = _RAND_4534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4535 = {1{`RANDOM}};
  _T_2457_im = _RAND_4535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4536 = {1{`RANDOM}};
  _T_2458_re = _RAND_4536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4537 = {1{`RANDOM}};
  _T_2458_im = _RAND_4537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4538 = {1{`RANDOM}};
  _T_2459_re = _RAND_4538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4539 = {1{`RANDOM}};
  _T_2459_im = _RAND_4539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4540 = {1{`RANDOM}};
  _T_2460_re = _RAND_4540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4541 = {1{`RANDOM}};
  _T_2460_im = _RAND_4541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4542 = {1{`RANDOM}};
  _T_2461_re = _RAND_4542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4543 = {1{`RANDOM}};
  _T_2461_im = _RAND_4543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4544 = {1{`RANDOM}};
  _T_2462_re = _RAND_4544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4545 = {1{`RANDOM}};
  _T_2462_im = _RAND_4545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4546 = {1{`RANDOM}};
  _T_2463_re = _RAND_4546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4547 = {1{`RANDOM}};
  _T_2463_im = _RAND_4547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4548 = {1{`RANDOM}};
  _T_2464_re = _RAND_4548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4549 = {1{`RANDOM}};
  _T_2464_im = _RAND_4549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4550 = {1{`RANDOM}};
  _T_2465_re = _RAND_4550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4551 = {1{`RANDOM}};
  _T_2465_im = _RAND_4551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4552 = {1{`RANDOM}};
  _T_2466_re = _RAND_4552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4553 = {1{`RANDOM}};
  _T_2466_im = _RAND_4553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4554 = {1{`RANDOM}};
  _T_2467_re = _RAND_4554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4555 = {1{`RANDOM}};
  _T_2467_im = _RAND_4555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4556 = {1{`RANDOM}};
  _T_2468_re = _RAND_4556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4557 = {1{`RANDOM}};
  _T_2468_im = _RAND_4557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4558 = {1{`RANDOM}};
  _T_2469_re = _RAND_4558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4559 = {1{`RANDOM}};
  _T_2469_im = _RAND_4559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4560 = {1{`RANDOM}};
  _T_2470_re = _RAND_4560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4561 = {1{`RANDOM}};
  _T_2470_im = _RAND_4561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4562 = {1{`RANDOM}};
  _T_2471_re = _RAND_4562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4563 = {1{`RANDOM}};
  _T_2471_im = _RAND_4563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4564 = {1{`RANDOM}};
  _T_2472_re = _RAND_4564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4565 = {1{`RANDOM}};
  _T_2472_im = _RAND_4565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4566 = {1{`RANDOM}};
  _T_2473_re = _RAND_4566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4567 = {1{`RANDOM}};
  _T_2473_im = _RAND_4567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4568 = {1{`RANDOM}};
  _T_2474_re = _RAND_4568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4569 = {1{`RANDOM}};
  _T_2474_im = _RAND_4569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4570 = {1{`RANDOM}};
  _T_2475_re = _RAND_4570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4571 = {1{`RANDOM}};
  _T_2475_im = _RAND_4571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4572 = {1{`RANDOM}};
  _T_2476_re = _RAND_4572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4573 = {1{`RANDOM}};
  _T_2476_im = _RAND_4573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4574 = {1{`RANDOM}};
  _T_2477_re = _RAND_4574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4575 = {1{`RANDOM}};
  _T_2477_im = _RAND_4575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4576 = {1{`RANDOM}};
  _T_2478_re = _RAND_4576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4577 = {1{`RANDOM}};
  _T_2478_im = _RAND_4577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4578 = {1{`RANDOM}};
  _T_2479_re = _RAND_4578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4579 = {1{`RANDOM}};
  _T_2479_im = _RAND_4579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4580 = {1{`RANDOM}};
  _T_2480_re = _RAND_4580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4581 = {1{`RANDOM}};
  _T_2480_im = _RAND_4581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4582 = {1{`RANDOM}};
  _T_2481_re = _RAND_4582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4583 = {1{`RANDOM}};
  _T_2481_im = _RAND_4583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4584 = {1{`RANDOM}};
  _T_2482_re = _RAND_4584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4585 = {1{`RANDOM}};
  _T_2482_im = _RAND_4585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4586 = {1{`RANDOM}};
  _T_2483_re = _RAND_4586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4587 = {1{`RANDOM}};
  _T_2483_im = _RAND_4587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4588 = {1{`RANDOM}};
  _T_2484_re = _RAND_4588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4589 = {1{`RANDOM}};
  _T_2484_im = _RAND_4589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4590 = {1{`RANDOM}};
  _T_2485_re = _RAND_4590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4591 = {1{`RANDOM}};
  _T_2485_im = _RAND_4591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4592 = {1{`RANDOM}};
  _T_2486_re = _RAND_4592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4593 = {1{`RANDOM}};
  _T_2486_im = _RAND_4593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4594 = {1{`RANDOM}};
  _T_2487_re = _RAND_4594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4595 = {1{`RANDOM}};
  _T_2487_im = _RAND_4595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4596 = {1{`RANDOM}};
  _T_2488_re = _RAND_4596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4597 = {1{`RANDOM}};
  _T_2488_im = _RAND_4597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4598 = {1{`RANDOM}};
  _T_2489_re = _RAND_4598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4599 = {1{`RANDOM}};
  _T_2489_im = _RAND_4599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4600 = {1{`RANDOM}};
  _T_2490_re = _RAND_4600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4601 = {1{`RANDOM}};
  _T_2490_im = _RAND_4601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4602 = {1{`RANDOM}};
  _T_2491_re = _RAND_4602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4603 = {1{`RANDOM}};
  _T_2491_im = _RAND_4603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4604 = {1{`RANDOM}};
  _T_2492_re = _RAND_4604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4605 = {1{`RANDOM}};
  _T_2492_im = _RAND_4605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4606 = {1{`RANDOM}};
  _T_2493_re = _RAND_4606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4607 = {1{`RANDOM}};
  _T_2493_im = _RAND_4607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4608 = {1{`RANDOM}};
  _T_2494_re = _RAND_4608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4609 = {1{`RANDOM}};
  _T_2494_im = _RAND_4609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4610 = {1{`RANDOM}};
  _T_2495_re = _RAND_4610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4611 = {1{`RANDOM}};
  _T_2495_im = _RAND_4611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4612 = {1{`RANDOM}};
  _T_2496_re = _RAND_4612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4613 = {1{`RANDOM}};
  _T_2496_im = _RAND_4613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4614 = {1{`RANDOM}};
  _T_2497_re = _RAND_4614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4615 = {1{`RANDOM}};
  _T_2497_im = _RAND_4615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4616 = {1{`RANDOM}};
  _T_2498_re = _RAND_4616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4617 = {1{`RANDOM}};
  _T_2498_im = _RAND_4617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4618 = {1{`RANDOM}};
  _T_2499_re = _RAND_4618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4619 = {1{`RANDOM}};
  _T_2499_im = _RAND_4619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4620 = {1{`RANDOM}};
  _T_2500_re = _RAND_4620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4621 = {1{`RANDOM}};
  _T_2500_im = _RAND_4621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4622 = {1{`RANDOM}};
  _T_2501_re = _RAND_4622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4623 = {1{`RANDOM}};
  _T_2501_im = _RAND_4623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4624 = {1{`RANDOM}};
  _T_2502_re = _RAND_4624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4625 = {1{`RANDOM}};
  _T_2502_im = _RAND_4625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4626 = {1{`RANDOM}};
  _T_2503_re = _RAND_4626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4627 = {1{`RANDOM}};
  _T_2503_im = _RAND_4627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4628 = {1{`RANDOM}};
  _T_2504_re = _RAND_4628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4629 = {1{`RANDOM}};
  _T_2504_im = _RAND_4629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4630 = {1{`RANDOM}};
  _T_2505_re = _RAND_4630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4631 = {1{`RANDOM}};
  _T_2505_im = _RAND_4631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4632 = {1{`RANDOM}};
  _T_2506_re = _RAND_4632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4633 = {1{`RANDOM}};
  _T_2506_im = _RAND_4633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4634 = {1{`RANDOM}};
  _T_2507_re = _RAND_4634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4635 = {1{`RANDOM}};
  _T_2507_im = _RAND_4635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4636 = {1{`RANDOM}};
  _T_2508_re = _RAND_4636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4637 = {1{`RANDOM}};
  _T_2508_im = _RAND_4637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4638 = {1{`RANDOM}};
  _T_2509_re = _RAND_4638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4639 = {1{`RANDOM}};
  _T_2509_im = _RAND_4639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4640 = {1{`RANDOM}};
  _T_2510_re = _RAND_4640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4641 = {1{`RANDOM}};
  _T_2510_im = _RAND_4641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4642 = {1{`RANDOM}};
  _T_2511_re = _RAND_4642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4643 = {1{`RANDOM}};
  _T_2511_im = _RAND_4643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4644 = {1{`RANDOM}};
  _T_2512_re = _RAND_4644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4645 = {1{`RANDOM}};
  _T_2512_im = _RAND_4645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4646 = {1{`RANDOM}};
  _T_2513_re = _RAND_4646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4647 = {1{`RANDOM}};
  _T_2513_im = _RAND_4647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4648 = {1{`RANDOM}};
  _T_2514_re = _RAND_4648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4649 = {1{`RANDOM}};
  _T_2514_im = _RAND_4649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4650 = {1{`RANDOM}};
  _T_2515_re = _RAND_4650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4651 = {1{`RANDOM}};
  _T_2515_im = _RAND_4651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4652 = {1{`RANDOM}};
  _T_2516_re = _RAND_4652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4653 = {1{`RANDOM}};
  _T_2516_im = _RAND_4653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4654 = {1{`RANDOM}};
  _T_2517_re = _RAND_4654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4655 = {1{`RANDOM}};
  _T_2517_im = _RAND_4655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4656 = {1{`RANDOM}};
  _T_2518_re = _RAND_4656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4657 = {1{`RANDOM}};
  _T_2518_im = _RAND_4657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4658 = {1{`RANDOM}};
  _T_2519_re = _RAND_4658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4659 = {1{`RANDOM}};
  _T_2519_im = _RAND_4659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4660 = {1{`RANDOM}};
  _T_2520_re = _RAND_4660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4661 = {1{`RANDOM}};
  _T_2520_im = _RAND_4661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4662 = {1{`RANDOM}};
  _T_2521_re = _RAND_4662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4663 = {1{`RANDOM}};
  _T_2521_im = _RAND_4663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4664 = {1{`RANDOM}};
  _T_2522_re = _RAND_4664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4665 = {1{`RANDOM}};
  _T_2522_im = _RAND_4665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4666 = {1{`RANDOM}};
  _T_2523_re = _RAND_4666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4667 = {1{`RANDOM}};
  _T_2523_im = _RAND_4667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4668 = {1{`RANDOM}};
  _T_2524_re = _RAND_4668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4669 = {1{`RANDOM}};
  _T_2524_im = _RAND_4669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4670 = {1{`RANDOM}};
  _T_2525_re = _RAND_4670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4671 = {1{`RANDOM}};
  _T_2525_im = _RAND_4671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4672 = {1{`RANDOM}};
  _T_2526_re = _RAND_4672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4673 = {1{`RANDOM}};
  _T_2526_im = _RAND_4673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4674 = {1{`RANDOM}};
  _T_2527_re = _RAND_4674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4675 = {1{`RANDOM}};
  _T_2527_im = _RAND_4675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4676 = {1{`RANDOM}};
  _T_2528_re = _RAND_4676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4677 = {1{`RANDOM}};
  _T_2528_im = _RAND_4677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4678 = {1{`RANDOM}};
  _T_2529_re = _RAND_4678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4679 = {1{`RANDOM}};
  _T_2529_im = _RAND_4679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4680 = {1{`RANDOM}};
  _T_2530_re = _RAND_4680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4681 = {1{`RANDOM}};
  _T_2530_im = _RAND_4681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4682 = {1{`RANDOM}};
  _T_2531_re = _RAND_4682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4683 = {1{`RANDOM}};
  _T_2531_im = _RAND_4683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4684 = {1{`RANDOM}};
  _T_2532_re = _RAND_4684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4685 = {1{`RANDOM}};
  _T_2532_im = _RAND_4685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4686 = {1{`RANDOM}};
  _T_2533_re = _RAND_4686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4687 = {1{`RANDOM}};
  _T_2533_im = _RAND_4687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4688 = {1{`RANDOM}};
  _T_2534_re = _RAND_4688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4689 = {1{`RANDOM}};
  _T_2534_im = _RAND_4689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4690 = {1{`RANDOM}};
  _T_2535_re = _RAND_4690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4691 = {1{`RANDOM}};
  _T_2535_im = _RAND_4691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4692 = {1{`RANDOM}};
  _T_2536_re = _RAND_4692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4693 = {1{`RANDOM}};
  _T_2536_im = _RAND_4693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4694 = {1{`RANDOM}};
  _T_2537_re = _RAND_4694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4695 = {1{`RANDOM}};
  _T_2537_im = _RAND_4695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4696 = {1{`RANDOM}};
  _T_2538_re = _RAND_4696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4697 = {1{`RANDOM}};
  _T_2538_im = _RAND_4697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4698 = {1{`RANDOM}};
  _T_2539_re = _RAND_4698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4699 = {1{`RANDOM}};
  _T_2539_im = _RAND_4699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4700 = {1{`RANDOM}};
  _T_2540_re = _RAND_4700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4701 = {1{`RANDOM}};
  _T_2540_im = _RAND_4701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4702 = {1{`RANDOM}};
  _T_2541_re = _RAND_4702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4703 = {1{`RANDOM}};
  _T_2541_im = _RAND_4703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4704 = {1{`RANDOM}};
  _T_2542_re = _RAND_4704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4705 = {1{`RANDOM}};
  _T_2542_im = _RAND_4705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4706 = {1{`RANDOM}};
  _T_2543_re = _RAND_4706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4707 = {1{`RANDOM}};
  _T_2543_im = _RAND_4707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4708 = {1{`RANDOM}};
  _T_2544_re = _RAND_4708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4709 = {1{`RANDOM}};
  _T_2544_im = _RAND_4709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4710 = {1{`RANDOM}};
  _T_2545_re = _RAND_4710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4711 = {1{`RANDOM}};
  _T_2545_im = _RAND_4711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4712 = {1{`RANDOM}};
  _T_2546_re = _RAND_4712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4713 = {1{`RANDOM}};
  _T_2546_im = _RAND_4713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4714 = {1{`RANDOM}};
  _T_2547_re = _RAND_4714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4715 = {1{`RANDOM}};
  _T_2547_im = _RAND_4715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4716 = {1{`RANDOM}};
  _T_2548_re = _RAND_4716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4717 = {1{`RANDOM}};
  _T_2548_im = _RAND_4717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4718 = {1{`RANDOM}};
  _T_2549_re = _RAND_4718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4719 = {1{`RANDOM}};
  _T_2549_im = _RAND_4719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4720 = {1{`RANDOM}};
  _T_2550_re = _RAND_4720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4721 = {1{`RANDOM}};
  _T_2550_im = _RAND_4721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4722 = {1{`RANDOM}};
  _T_2551_re = _RAND_4722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4723 = {1{`RANDOM}};
  _T_2551_im = _RAND_4723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4724 = {1{`RANDOM}};
  _T_2552_re = _RAND_4724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4725 = {1{`RANDOM}};
  _T_2552_im = _RAND_4725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4726 = {1{`RANDOM}};
  _T_2553_re = _RAND_4726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4727 = {1{`RANDOM}};
  _T_2553_im = _RAND_4727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4728 = {1{`RANDOM}};
  _T_2554_re = _RAND_4728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4729 = {1{`RANDOM}};
  _T_2554_im = _RAND_4729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4730 = {1{`RANDOM}};
  _T_2555_re = _RAND_4730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4731 = {1{`RANDOM}};
  _T_2555_im = _RAND_4731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4732 = {1{`RANDOM}};
  _T_2556_re = _RAND_4732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4733 = {1{`RANDOM}};
  _T_2556_im = _RAND_4733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4734 = {1{`RANDOM}};
  _T_2557_re = _RAND_4734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4735 = {1{`RANDOM}};
  _T_2557_im = _RAND_4735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4736 = {1{`RANDOM}};
  _T_2558_re = _RAND_4736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4737 = {1{`RANDOM}};
  _T_2558_im = _RAND_4737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4738 = {1{`RANDOM}};
  _T_2559_re = _RAND_4738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4739 = {1{`RANDOM}};
  _T_2559_im = _RAND_4739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4740 = {1{`RANDOM}};
  _T_2560_re = _RAND_4740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4741 = {1{`RANDOM}};
  _T_2560_im = _RAND_4741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4742 = {1{`RANDOM}};
  _T_2561_re = _RAND_4742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4743 = {1{`RANDOM}};
  _T_2561_im = _RAND_4743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4744 = {1{`RANDOM}};
  _T_2562_re = _RAND_4744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4745 = {1{`RANDOM}};
  _T_2562_im = _RAND_4745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4746 = {1{`RANDOM}};
  _T_2563_re = _RAND_4746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4747 = {1{`RANDOM}};
  _T_2563_im = _RAND_4747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4748 = {1{`RANDOM}};
  _T_2564_re = _RAND_4748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4749 = {1{`RANDOM}};
  _T_2564_im = _RAND_4749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4750 = {1{`RANDOM}};
  _T_2565_re = _RAND_4750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4751 = {1{`RANDOM}};
  _T_2565_im = _RAND_4751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4752 = {1{`RANDOM}};
  _T_2566_re = _RAND_4752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4753 = {1{`RANDOM}};
  _T_2566_im = _RAND_4753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4754 = {1{`RANDOM}};
  _T_2567_re = _RAND_4754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4755 = {1{`RANDOM}};
  _T_2567_im = _RAND_4755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4756 = {1{`RANDOM}};
  _T_2568_re = _RAND_4756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4757 = {1{`RANDOM}};
  _T_2568_im = _RAND_4757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4758 = {1{`RANDOM}};
  _T_2569_re = _RAND_4758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4759 = {1{`RANDOM}};
  _T_2569_im = _RAND_4759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4760 = {1{`RANDOM}};
  _T_2570_re = _RAND_4760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4761 = {1{`RANDOM}};
  _T_2570_im = _RAND_4761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4762 = {1{`RANDOM}};
  _T_2571_re = _RAND_4762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4763 = {1{`RANDOM}};
  _T_2571_im = _RAND_4763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4764 = {1{`RANDOM}};
  _T_2572_re = _RAND_4764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4765 = {1{`RANDOM}};
  _T_2572_im = _RAND_4765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4766 = {1{`RANDOM}};
  _T_2573_re = _RAND_4766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4767 = {1{`RANDOM}};
  _T_2573_im = _RAND_4767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4768 = {1{`RANDOM}};
  _T_2574_re = _RAND_4768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4769 = {1{`RANDOM}};
  _T_2574_im = _RAND_4769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4770 = {1{`RANDOM}};
  _T_2575_re = _RAND_4770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4771 = {1{`RANDOM}};
  _T_2575_im = _RAND_4771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4772 = {1{`RANDOM}};
  _T_2576_re = _RAND_4772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4773 = {1{`RANDOM}};
  _T_2576_im = _RAND_4773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4774 = {1{`RANDOM}};
  _T_2577_re = _RAND_4774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4775 = {1{`RANDOM}};
  _T_2577_im = _RAND_4775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4776 = {1{`RANDOM}};
  _T_2578_re = _RAND_4776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4777 = {1{`RANDOM}};
  _T_2578_im = _RAND_4777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4778 = {1{`RANDOM}};
  _T_2579_re = _RAND_4778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4779 = {1{`RANDOM}};
  _T_2579_im = _RAND_4779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4780 = {1{`RANDOM}};
  _T_2580_re = _RAND_4780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4781 = {1{`RANDOM}};
  _T_2580_im = _RAND_4781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4782 = {1{`RANDOM}};
  _T_2581_re = _RAND_4782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4783 = {1{`RANDOM}};
  _T_2581_im = _RAND_4783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4784 = {1{`RANDOM}};
  _T_2582_re = _RAND_4784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4785 = {1{`RANDOM}};
  _T_2582_im = _RAND_4785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4786 = {1{`RANDOM}};
  _T_2583_re = _RAND_4786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4787 = {1{`RANDOM}};
  _T_2583_im = _RAND_4787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4788 = {1{`RANDOM}};
  _T_2584_re = _RAND_4788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4789 = {1{`RANDOM}};
  _T_2584_im = _RAND_4789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4790 = {1{`RANDOM}};
  _T_2585_re = _RAND_4790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4791 = {1{`RANDOM}};
  _T_2585_im = _RAND_4791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4792 = {1{`RANDOM}};
  _T_2586_re = _RAND_4792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4793 = {1{`RANDOM}};
  _T_2586_im = _RAND_4793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4794 = {1{`RANDOM}};
  _T_2587_re = _RAND_4794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4795 = {1{`RANDOM}};
  _T_2587_im = _RAND_4795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4796 = {1{`RANDOM}};
  _T_2588_re = _RAND_4796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4797 = {1{`RANDOM}};
  _T_2588_im = _RAND_4797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4798 = {1{`RANDOM}};
  _T_2589_re = _RAND_4798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4799 = {1{`RANDOM}};
  _T_2589_im = _RAND_4799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4800 = {1{`RANDOM}};
  _T_2590_re = _RAND_4800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4801 = {1{`RANDOM}};
  _T_2590_im = _RAND_4801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4802 = {1{`RANDOM}};
  _T_2591_re = _RAND_4802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4803 = {1{`RANDOM}};
  _T_2591_im = _RAND_4803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4804 = {1{`RANDOM}};
  _T_2592_re = _RAND_4804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4805 = {1{`RANDOM}};
  _T_2592_im = _RAND_4805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4806 = {1{`RANDOM}};
  _T_2593_re = _RAND_4806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4807 = {1{`RANDOM}};
  _T_2593_im = _RAND_4807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4808 = {1{`RANDOM}};
  _T_2594_re = _RAND_4808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4809 = {1{`RANDOM}};
  _T_2594_im = _RAND_4809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4810 = {1{`RANDOM}};
  _T_2595_re = _RAND_4810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4811 = {1{`RANDOM}};
  _T_2595_im = _RAND_4811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4812 = {1{`RANDOM}};
  _T_2596_re = _RAND_4812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4813 = {1{`RANDOM}};
  _T_2596_im = _RAND_4813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4814 = {1{`RANDOM}};
  _T_2597_re = _RAND_4814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4815 = {1{`RANDOM}};
  _T_2597_im = _RAND_4815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4816 = {1{`RANDOM}};
  _T_2598_re = _RAND_4816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4817 = {1{`RANDOM}};
  _T_2598_im = _RAND_4817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4818 = {1{`RANDOM}};
  _T_2599_re = _RAND_4818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4819 = {1{`RANDOM}};
  _T_2599_im = _RAND_4819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4820 = {1{`RANDOM}};
  _T_2600_re = _RAND_4820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4821 = {1{`RANDOM}};
  _T_2600_im = _RAND_4821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4822 = {1{`RANDOM}};
  _T_2601_re = _RAND_4822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4823 = {1{`RANDOM}};
  _T_2601_im = _RAND_4823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4824 = {1{`RANDOM}};
  _T_2602_re = _RAND_4824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4825 = {1{`RANDOM}};
  _T_2602_im = _RAND_4825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4826 = {1{`RANDOM}};
  _T_2603_re = _RAND_4826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4827 = {1{`RANDOM}};
  _T_2603_im = _RAND_4827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4828 = {1{`RANDOM}};
  _T_2604_re = _RAND_4828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4829 = {1{`RANDOM}};
  _T_2604_im = _RAND_4829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4830 = {1{`RANDOM}};
  _T_2605_re = _RAND_4830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4831 = {1{`RANDOM}};
  _T_2605_im = _RAND_4831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4832 = {1{`RANDOM}};
  _T_2606_re = _RAND_4832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4833 = {1{`RANDOM}};
  _T_2606_im = _RAND_4833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4834 = {1{`RANDOM}};
  _T_2607_re = _RAND_4834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4835 = {1{`RANDOM}};
  _T_2607_im = _RAND_4835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4836 = {1{`RANDOM}};
  _T_2608_re = _RAND_4836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4837 = {1{`RANDOM}};
  _T_2608_im = _RAND_4837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4838 = {1{`RANDOM}};
  _T_2609_re = _RAND_4838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4839 = {1{`RANDOM}};
  _T_2609_im = _RAND_4839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4840 = {1{`RANDOM}};
  _T_2610_re = _RAND_4840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4841 = {1{`RANDOM}};
  _T_2610_im = _RAND_4841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4842 = {1{`RANDOM}};
  _T_2611_re = _RAND_4842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4843 = {1{`RANDOM}};
  _T_2611_im = _RAND_4843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4844 = {1{`RANDOM}};
  _T_2612_re = _RAND_4844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4845 = {1{`RANDOM}};
  _T_2612_im = _RAND_4845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4846 = {1{`RANDOM}};
  _T_2613_re = _RAND_4846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4847 = {1{`RANDOM}};
  _T_2613_im = _RAND_4847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4848 = {1{`RANDOM}};
  _T_2614_re = _RAND_4848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4849 = {1{`RANDOM}};
  _T_2614_im = _RAND_4849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4850 = {1{`RANDOM}};
  _T_2615_re = _RAND_4850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4851 = {1{`RANDOM}};
  _T_2615_im = _RAND_4851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4852 = {1{`RANDOM}};
  _T_2616_re = _RAND_4852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4853 = {1{`RANDOM}};
  _T_2616_im = _RAND_4853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4854 = {1{`RANDOM}};
  _T_2617_re = _RAND_4854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4855 = {1{`RANDOM}};
  _T_2617_im = _RAND_4855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4856 = {1{`RANDOM}};
  _T_2618_re = _RAND_4856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4857 = {1{`RANDOM}};
  _T_2618_im = _RAND_4857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4858 = {1{`RANDOM}};
  _T_2619_re = _RAND_4858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4859 = {1{`RANDOM}};
  _T_2619_im = _RAND_4859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4860 = {1{`RANDOM}};
  _T_2620_re = _RAND_4860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4861 = {1{`RANDOM}};
  _T_2620_im = _RAND_4861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4862 = {1{`RANDOM}};
  _T_2621_re = _RAND_4862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4863 = {1{`RANDOM}};
  _T_2621_im = _RAND_4863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4864 = {1{`RANDOM}};
  _T_2622_re = _RAND_4864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4865 = {1{`RANDOM}};
  _T_2622_im = _RAND_4865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4866 = {1{`RANDOM}};
  _T_2623_re = _RAND_4866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4867 = {1{`RANDOM}};
  _T_2623_im = _RAND_4867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4868 = {1{`RANDOM}};
  _T_2624_re = _RAND_4868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4869 = {1{`RANDOM}};
  _T_2624_im = _RAND_4869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4870 = {1{`RANDOM}};
  _T_2625_re = _RAND_4870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4871 = {1{`RANDOM}};
  _T_2625_im = _RAND_4871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4872 = {1{`RANDOM}};
  _T_2626_re = _RAND_4872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4873 = {1{`RANDOM}};
  _T_2626_im = _RAND_4873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4874 = {1{`RANDOM}};
  _T_2627_re = _RAND_4874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4875 = {1{`RANDOM}};
  _T_2627_im = _RAND_4875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4876 = {1{`RANDOM}};
  _T_2628_re = _RAND_4876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4877 = {1{`RANDOM}};
  _T_2628_im = _RAND_4877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4878 = {1{`RANDOM}};
  _T_2629_re = _RAND_4878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4879 = {1{`RANDOM}};
  _T_2629_im = _RAND_4879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4880 = {1{`RANDOM}};
  _T_2630_re = _RAND_4880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4881 = {1{`RANDOM}};
  _T_2630_im = _RAND_4881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4882 = {1{`RANDOM}};
  _T_2631_re = _RAND_4882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4883 = {1{`RANDOM}};
  _T_2631_im = _RAND_4883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4884 = {1{`RANDOM}};
  _T_2632_re = _RAND_4884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4885 = {1{`RANDOM}};
  _T_2632_im = _RAND_4885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4886 = {1{`RANDOM}};
  _T_2633_re = _RAND_4886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4887 = {1{`RANDOM}};
  _T_2633_im = _RAND_4887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4888 = {1{`RANDOM}};
  _T_2634_re = _RAND_4888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4889 = {1{`RANDOM}};
  _T_2634_im = _RAND_4889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4890 = {1{`RANDOM}};
  _T_2635_re = _RAND_4890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4891 = {1{`RANDOM}};
  _T_2635_im = _RAND_4891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4892 = {1{`RANDOM}};
  _T_2636_re = _RAND_4892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4893 = {1{`RANDOM}};
  _T_2636_im = _RAND_4893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4894 = {1{`RANDOM}};
  _T_2637_re = _RAND_4894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4895 = {1{`RANDOM}};
  _T_2637_im = _RAND_4895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4896 = {1{`RANDOM}};
  _T_2638_re = _RAND_4896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4897 = {1{`RANDOM}};
  _T_2638_im = _RAND_4897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4898 = {1{`RANDOM}};
  _T_2639_re = _RAND_4898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4899 = {1{`RANDOM}};
  _T_2639_im = _RAND_4899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4900 = {1{`RANDOM}};
  _T_2640_re = _RAND_4900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4901 = {1{`RANDOM}};
  _T_2640_im = _RAND_4901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4902 = {1{`RANDOM}};
  _T_2641_re = _RAND_4902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4903 = {1{`RANDOM}};
  _T_2641_im = _RAND_4903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4904 = {1{`RANDOM}};
  _T_2642_re = _RAND_4904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4905 = {1{`RANDOM}};
  _T_2642_im = _RAND_4905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4906 = {1{`RANDOM}};
  _T_2643_re = _RAND_4906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4907 = {1{`RANDOM}};
  _T_2643_im = _RAND_4907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4908 = {1{`RANDOM}};
  _T_2644_re = _RAND_4908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4909 = {1{`RANDOM}};
  _T_2644_im = _RAND_4909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4910 = {1{`RANDOM}};
  _T_2645_re = _RAND_4910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4911 = {1{`RANDOM}};
  _T_2645_im = _RAND_4911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4912 = {1{`RANDOM}};
  _T_2646_re = _RAND_4912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4913 = {1{`RANDOM}};
  _T_2646_im = _RAND_4913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4914 = {1{`RANDOM}};
  _T_2647_re = _RAND_4914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4915 = {1{`RANDOM}};
  _T_2647_im = _RAND_4915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4916 = {1{`RANDOM}};
  _T_2648_re = _RAND_4916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4917 = {1{`RANDOM}};
  _T_2648_im = _RAND_4917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4918 = {1{`RANDOM}};
  _T_2649_re = _RAND_4918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4919 = {1{`RANDOM}};
  _T_2649_im = _RAND_4919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4920 = {1{`RANDOM}};
  _T_2650_re = _RAND_4920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4921 = {1{`RANDOM}};
  _T_2650_im = _RAND_4921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4922 = {1{`RANDOM}};
  _T_2651_re = _RAND_4922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4923 = {1{`RANDOM}};
  _T_2651_im = _RAND_4923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4924 = {1{`RANDOM}};
  _T_2652_re = _RAND_4924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4925 = {1{`RANDOM}};
  _T_2652_im = _RAND_4925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4926 = {1{`RANDOM}};
  _T_2653_re = _RAND_4926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4927 = {1{`RANDOM}};
  _T_2653_im = _RAND_4927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4928 = {1{`RANDOM}};
  _T_2654_re = _RAND_4928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4929 = {1{`RANDOM}};
  _T_2654_im = _RAND_4929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4930 = {1{`RANDOM}};
  _T_2655_re = _RAND_4930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4931 = {1{`RANDOM}};
  _T_2655_im = _RAND_4931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4932 = {1{`RANDOM}};
  _T_2656_re = _RAND_4932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4933 = {1{`RANDOM}};
  _T_2656_im = _RAND_4933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4934 = {1{`RANDOM}};
  _T_2657_re = _RAND_4934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4935 = {1{`RANDOM}};
  _T_2657_im = _RAND_4935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4936 = {1{`RANDOM}};
  _T_2658_re = _RAND_4936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4937 = {1{`RANDOM}};
  _T_2658_im = _RAND_4937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4938 = {1{`RANDOM}};
  _T_2659_re = _RAND_4938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4939 = {1{`RANDOM}};
  _T_2659_im = _RAND_4939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4940 = {1{`RANDOM}};
  _T_2660_re = _RAND_4940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4941 = {1{`RANDOM}};
  _T_2660_im = _RAND_4941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4942 = {1{`RANDOM}};
  _T_2661_re = _RAND_4942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4943 = {1{`RANDOM}};
  _T_2661_im = _RAND_4943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4944 = {1{`RANDOM}};
  _T_2662_re = _RAND_4944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4945 = {1{`RANDOM}};
  _T_2662_im = _RAND_4945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4946 = {1{`RANDOM}};
  _T_2663_re = _RAND_4946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4947 = {1{`RANDOM}};
  _T_2663_im = _RAND_4947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4948 = {1{`RANDOM}};
  _T_2664_re = _RAND_4948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4949 = {1{`RANDOM}};
  _T_2664_im = _RAND_4949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4950 = {1{`RANDOM}};
  _T_2665_re = _RAND_4950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4951 = {1{`RANDOM}};
  _T_2665_im = _RAND_4951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4952 = {1{`RANDOM}};
  _T_2666_re = _RAND_4952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4953 = {1{`RANDOM}};
  _T_2666_im = _RAND_4953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4954 = {1{`RANDOM}};
  _T_2667_re = _RAND_4954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4955 = {1{`RANDOM}};
  _T_2667_im = _RAND_4955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4956 = {1{`RANDOM}};
  _T_2668_re = _RAND_4956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4957 = {1{`RANDOM}};
  _T_2668_im = _RAND_4957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4958 = {1{`RANDOM}};
  _T_2669_re = _RAND_4958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4959 = {1{`RANDOM}};
  _T_2669_im = _RAND_4959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4960 = {1{`RANDOM}};
  _T_2670_re = _RAND_4960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4961 = {1{`RANDOM}};
  _T_2670_im = _RAND_4961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4962 = {1{`RANDOM}};
  _T_2671_re = _RAND_4962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4963 = {1{`RANDOM}};
  _T_2671_im = _RAND_4963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4964 = {1{`RANDOM}};
  _T_2672_re = _RAND_4964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4965 = {1{`RANDOM}};
  _T_2672_im = _RAND_4965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4966 = {1{`RANDOM}};
  _T_2673_re = _RAND_4966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4967 = {1{`RANDOM}};
  _T_2673_im = _RAND_4967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4968 = {1{`RANDOM}};
  _T_2674_re = _RAND_4968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4969 = {1{`RANDOM}};
  _T_2674_im = _RAND_4969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4970 = {1{`RANDOM}};
  _T_2675_re = _RAND_4970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4971 = {1{`RANDOM}};
  _T_2675_im = _RAND_4971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4972 = {1{`RANDOM}};
  _T_2676_re = _RAND_4972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4973 = {1{`RANDOM}};
  _T_2676_im = _RAND_4973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4974 = {1{`RANDOM}};
  _T_2677_re = _RAND_4974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4975 = {1{`RANDOM}};
  _T_2677_im = _RAND_4975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4976 = {1{`RANDOM}};
  _T_2678_re = _RAND_4976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4977 = {1{`RANDOM}};
  _T_2678_im = _RAND_4977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4978 = {1{`RANDOM}};
  _T_2679_re = _RAND_4978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4979 = {1{`RANDOM}};
  _T_2679_im = _RAND_4979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4980 = {1{`RANDOM}};
  _T_2680_re = _RAND_4980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4981 = {1{`RANDOM}};
  _T_2680_im = _RAND_4981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4982 = {1{`RANDOM}};
  _T_2681_re = _RAND_4982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4983 = {1{`RANDOM}};
  _T_2681_im = _RAND_4983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4984 = {1{`RANDOM}};
  _T_2682_re = _RAND_4984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4985 = {1{`RANDOM}};
  _T_2682_im = _RAND_4985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4986 = {1{`RANDOM}};
  _T_2683_re = _RAND_4986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4987 = {1{`RANDOM}};
  _T_2683_im = _RAND_4987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4988 = {1{`RANDOM}};
  _T_2684_re = _RAND_4988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4989 = {1{`RANDOM}};
  _T_2684_im = _RAND_4989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4990 = {1{`RANDOM}};
  _T_2685_re = _RAND_4990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4991 = {1{`RANDOM}};
  _T_2685_im = _RAND_4991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4992 = {1{`RANDOM}};
  _T_2686_re = _RAND_4992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4993 = {1{`RANDOM}};
  _T_2686_im = _RAND_4993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4994 = {1{`RANDOM}};
  _T_2687_re = _RAND_4994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4995 = {1{`RANDOM}};
  _T_2687_im = _RAND_4995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4996 = {1{`RANDOM}};
  _T_2688_re = _RAND_4996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4997 = {1{`RANDOM}};
  _T_2688_im = _RAND_4997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4998 = {1{`RANDOM}};
  _T_2689_re = _RAND_4998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4999 = {1{`RANDOM}};
  _T_2689_im = _RAND_4999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5000 = {1{`RANDOM}};
  _T_2690_re = _RAND_5000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5001 = {1{`RANDOM}};
  _T_2690_im = _RAND_5001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5002 = {1{`RANDOM}};
  _T_2691_re = _RAND_5002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5003 = {1{`RANDOM}};
  _T_2691_im = _RAND_5003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5004 = {1{`RANDOM}};
  _T_2692_re = _RAND_5004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5005 = {1{`RANDOM}};
  _T_2692_im = _RAND_5005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5006 = {1{`RANDOM}};
  _T_2693_re = _RAND_5006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5007 = {1{`RANDOM}};
  _T_2693_im = _RAND_5007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5008 = {1{`RANDOM}};
  _T_2694_re = _RAND_5008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5009 = {1{`RANDOM}};
  _T_2694_im = _RAND_5009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5010 = {1{`RANDOM}};
  _T_2695_re = _RAND_5010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5011 = {1{`RANDOM}};
  _T_2695_im = _RAND_5011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5012 = {1{`RANDOM}};
  _T_2696_re = _RAND_5012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5013 = {1{`RANDOM}};
  _T_2696_im = _RAND_5013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5014 = {1{`RANDOM}};
  _T_2697_re = _RAND_5014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5015 = {1{`RANDOM}};
  _T_2697_im = _RAND_5015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5016 = {1{`RANDOM}};
  _T_2698_re = _RAND_5016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5017 = {1{`RANDOM}};
  _T_2698_im = _RAND_5017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5018 = {1{`RANDOM}};
  _T_2699_re = _RAND_5018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5019 = {1{`RANDOM}};
  _T_2699_im = _RAND_5019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5020 = {1{`RANDOM}};
  _T_2700_re = _RAND_5020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5021 = {1{`RANDOM}};
  _T_2700_im = _RAND_5021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5022 = {1{`RANDOM}};
  _T_2701_re = _RAND_5022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5023 = {1{`RANDOM}};
  _T_2701_im = _RAND_5023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5024 = {1{`RANDOM}};
  _T_2702_re = _RAND_5024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5025 = {1{`RANDOM}};
  _T_2702_im = _RAND_5025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5026 = {1{`RANDOM}};
  _T_2703_re = _RAND_5026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5027 = {1{`RANDOM}};
  _T_2703_im = _RAND_5027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5028 = {1{`RANDOM}};
  _T_2704_re = _RAND_5028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5029 = {1{`RANDOM}};
  _T_2704_im = _RAND_5029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5030 = {1{`RANDOM}};
  _T_2705_re = _RAND_5030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5031 = {1{`RANDOM}};
  _T_2705_im = _RAND_5031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5032 = {1{`RANDOM}};
  _T_2706_re = _RAND_5032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5033 = {1{`RANDOM}};
  _T_2706_im = _RAND_5033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5034 = {1{`RANDOM}};
  _T_2707_re = _RAND_5034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5035 = {1{`RANDOM}};
  _T_2707_im = _RAND_5035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5036 = {1{`RANDOM}};
  _T_2708_re = _RAND_5036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5037 = {1{`RANDOM}};
  _T_2708_im = _RAND_5037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5038 = {1{`RANDOM}};
  _T_2709_re = _RAND_5038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5039 = {1{`RANDOM}};
  _T_2709_im = _RAND_5039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5040 = {1{`RANDOM}};
  _T_2710_re = _RAND_5040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5041 = {1{`RANDOM}};
  _T_2710_im = _RAND_5041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5042 = {1{`RANDOM}};
  _T_2711_re = _RAND_5042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5043 = {1{`RANDOM}};
  _T_2711_im = _RAND_5043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5044 = {1{`RANDOM}};
  _T_2712_re = _RAND_5044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5045 = {1{`RANDOM}};
  _T_2712_im = _RAND_5045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5046 = {1{`RANDOM}};
  _T_2713_re = _RAND_5046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5047 = {1{`RANDOM}};
  _T_2713_im = _RAND_5047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5048 = {1{`RANDOM}};
  _T_2714_re = _RAND_5048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5049 = {1{`RANDOM}};
  _T_2714_im = _RAND_5049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5050 = {1{`RANDOM}};
  _T_2715_re = _RAND_5050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5051 = {1{`RANDOM}};
  _T_2715_im = _RAND_5051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5052 = {1{`RANDOM}};
  _T_2716_re = _RAND_5052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5053 = {1{`RANDOM}};
  _T_2716_im = _RAND_5053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5054 = {1{`RANDOM}};
  _T_2717_re = _RAND_5054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5055 = {1{`RANDOM}};
  _T_2717_im = _RAND_5055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5056 = {1{`RANDOM}};
  _T_2718_re = _RAND_5056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5057 = {1{`RANDOM}};
  _T_2718_im = _RAND_5057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5058 = {1{`RANDOM}};
  _T_2719_re = _RAND_5058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5059 = {1{`RANDOM}};
  _T_2719_im = _RAND_5059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5060 = {1{`RANDOM}};
  _T_2720_re = _RAND_5060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5061 = {1{`RANDOM}};
  _T_2720_im = _RAND_5061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5062 = {1{`RANDOM}};
  _T_2721_re = _RAND_5062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5063 = {1{`RANDOM}};
  _T_2721_im = _RAND_5063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5064 = {1{`RANDOM}};
  _T_2722_re = _RAND_5064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5065 = {1{`RANDOM}};
  _T_2722_im = _RAND_5065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5066 = {1{`RANDOM}};
  _T_2723_re = _RAND_5066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5067 = {1{`RANDOM}};
  _T_2723_im = _RAND_5067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5068 = {1{`RANDOM}};
  _T_2724_re = _RAND_5068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5069 = {1{`RANDOM}};
  _T_2724_im = _RAND_5069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5070 = {1{`RANDOM}};
  _T_2725_re = _RAND_5070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5071 = {1{`RANDOM}};
  _T_2725_im = _RAND_5071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5072 = {1{`RANDOM}};
  _T_2726_re = _RAND_5072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5073 = {1{`RANDOM}};
  _T_2726_im = _RAND_5073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5074 = {1{`RANDOM}};
  _T_2727_re = _RAND_5074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5075 = {1{`RANDOM}};
  _T_2727_im = _RAND_5075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5076 = {1{`RANDOM}};
  _T_2728_re = _RAND_5076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5077 = {1{`RANDOM}};
  _T_2728_im = _RAND_5077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5078 = {1{`RANDOM}};
  _T_2729_re = _RAND_5078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5079 = {1{`RANDOM}};
  _T_2729_im = _RAND_5079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5080 = {1{`RANDOM}};
  _T_2730_re = _RAND_5080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5081 = {1{`RANDOM}};
  _T_2730_im = _RAND_5081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5082 = {1{`RANDOM}};
  _T_2731_re = _RAND_5082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5083 = {1{`RANDOM}};
  _T_2731_im = _RAND_5083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5084 = {1{`RANDOM}};
  _T_2732_re = _RAND_5084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5085 = {1{`RANDOM}};
  _T_2732_im = _RAND_5085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5086 = {1{`RANDOM}};
  _T_2733_re = _RAND_5086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5087 = {1{`RANDOM}};
  _T_2733_im = _RAND_5087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5088 = {1{`RANDOM}};
  _T_2734_re = _RAND_5088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5089 = {1{`RANDOM}};
  _T_2734_im = _RAND_5089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5090 = {1{`RANDOM}};
  _T_2735_re = _RAND_5090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5091 = {1{`RANDOM}};
  _T_2735_im = _RAND_5091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5092 = {1{`RANDOM}};
  _T_2736_re = _RAND_5092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5093 = {1{`RANDOM}};
  _T_2736_im = _RAND_5093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5094 = {1{`RANDOM}};
  _T_2737_re = _RAND_5094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5095 = {1{`RANDOM}};
  _T_2737_im = _RAND_5095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5096 = {1{`RANDOM}};
  _T_2738_re = _RAND_5096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5097 = {1{`RANDOM}};
  _T_2738_im = _RAND_5097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5098 = {1{`RANDOM}};
  _T_2739_re = _RAND_5098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5099 = {1{`RANDOM}};
  _T_2739_im = _RAND_5099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5100 = {1{`RANDOM}};
  _T_2740_re = _RAND_5100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5101 = {1{`RANDOM}};
  _T_2740_im = _RAND_5101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5102 = {1{`RANDOM}};
  _T_2741_re = _RAND_5102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5103 = {1{`RANDOM}};
  _T_2741_im = _RAND_5103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5104 = {1{`RANDOM}};
  _T_2742_re = _RAND_5104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5105 = {1{`RANDOM}};
  _T_2742_im = _RAND_5105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5106 = {1{`RANDOM}};
  _T_2743_re = _RAND_5106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5107 = {1{`RANDOM}};
  _T_2743_im = _RAND_5107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5108 = {1{`RANDOM}};
  _T_2744_re = _RAND_5108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5109 = {1{`RANDOM}};
  _T_2744_im = _RAND_5109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5110 = {1{`RANDOM}};
  _T_2745_re = _RAND_5110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5111 = {1{`RANDOM}};
  _T_2745_im = _RAND_5111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5112 = {1{`RANDOM}};
  _T_2746_re = _RAND_5112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5113 = {1{`RANDOM}};
  _T_2746_im = _RAND_5113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5114 = {1{`RANDOM}};
  _T_2747_re = _RAND_5114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5115 = {1{`RANDOM}};
  _T_2747_im = _RAND_5115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5116 = {1{`RANDOM}};
  _T_2748_re = _RAND_5116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5117 = {1{`RANDOM}};
  _T_2748_im = _RAND_5117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5118 = {1{`RANDOM}};
  _T_2749_re = _RAND_5118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5119 = {1{`RANDOM}};
  _T_2749_im = _RAND_5119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5120 = {1{`RANDOM}};
  _T_2750_re = _RAND_5120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5121 = {1{`RANDOM}};
  _T_2750_im = _RAND_5121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5122 = {1{`RANDOM}};
  _T_2751_re = _RAND_5122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5123 = {1{`RANDOM}};
  _T_2751_im = _RAND_5123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5124 = {1{`RANDOM}};
  _T_2752_re = _RAND_5124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5125 = {1{`RANDOM}};
  _T_2752_im = _RAND_5125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5126 = {1{`RANDOM}};
  _T_2753_re = _RAND_5126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5127 = {1{`RANDOM}};
  _T_2753_im = _RAND_5127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5128 = {1{`RANDOM}};
  _T_2754_re = _RAND_5128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5129 = {1{`RANDOM}};
  _T_2754_im = _RAND_5129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5130 = {1{`RANDOM}};
  _T_2755_re = _RAND_5130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5131 = {1{`RANDOM}};
  _T_2755_im = _RAND_5131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5132 = {1{`RANDOM}};
  _T_2756_re = _RAND_5132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5133 = {1{`RANDOM}};
  _T_2756_im = _RAND_5133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5134 = {1{`RANDOM}};
  _T_2757_re = _RAND_5134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5135 = {1{`RANDOM}};
  _T_2757_im = _RAND_5135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5136 = {1{`RANDOM}};
  _T_2758_re = _RAND_5136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5137 = {1{`RANDOM}};
  _T_2758_im = _RAND_5137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5138 = {1{`RANDOM}};
  _T_2759_re = _RAND_5138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5139 = {1{`RANDOM}};
  _T_2759_im = _RAND_5139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5140 = {1{`RANDOM}};
  _T_2760_re = _RAND_5140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5141 = {1{`RANDOM}};
  _T_2760_im = _RAND_5141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5142 = {1{`RANDOM}};
  _T_2761_re = _RAND_5142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5143 = {1{`RANDOM}};
  _T_2761_im = _RAND_5143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5144 = {1{`RANDOM}};
  _T_2762_re = _RAND_5144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5145 = {1{`RANDOM}};
  _T_2762_im = _RAND_5145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5146 = {1{`RANDOM}};
  _T_2763_re = _RAND_5146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5147 = {1{`RANDOM}};
  _T_2763_im = _RAND_5147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5148 = {1{`RANDOM}};
  _T_2764_re = _RAND_5148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5149 = {1{`RANDOM}};
  _T_2764_im = _RAND_5149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5150 = {1{`RANDOM}};
  _T_2765_re = _RAND_5150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5151 = {1{`RANDOM}};
  _T_2765_im = _RAND_5151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5152 = {1{`RANDOM}};
  _T_2766_re = _RAND_5152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5153 = {1{`RANDOM}};
  _T_2766_im = _RAND_5153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5154 = {1{`RANDOM}};
  _T_2767_re = _RAND_5154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5155 = {1{`RANDOM}};
  _T_2767_im = _RAND_5155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5156 = {1{`RANDOM}};
  _T_2768_re = _RAND_5156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5157 = {1{`RANDOM}};
  _T_2768_im = _RAND_5157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5158 = {1{`RANDOM}};
  _T_2769_re = _RAND_5158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5159 = {1{`RANDOM}};
  _T_2769_im = _RAND_5159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5160 = {1{`RANDOM}};
  _T_2770_re = _RAND_5160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5161 = {1{`RANDOM}};
  _T_2770_im = _RAND_5161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5162 = {1{`RANDOM}};
  _T_2771_re = _RAND_5162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5163 = {1{`RANDOM}};
  _T_2771_im = _RAND_5163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5164 = {1{`RANDOM}};
  _T_2772_re = _RAND_5164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5165 = {1{`RANDOM}};
  _T_2772_im = _RAND_5165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5166 = {1{`RANDOM}};
  _T_2773_re = _RAND_5166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5167 = {1{`RANDOM}};
  _T_2773_im = _RAND_5167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5168 = {1{`RANDOM}};
  _T_2774_re = _RAND_5168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5169 = {1{`RANDOM}};
  _T_2774_im = _RAND_5169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5170 = {1{`RANDOM}};
  _T_2775_re = _RAND_5170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5171 = {1{`RANDOM}};
  _T_2775_im = _RAND_5171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5172 = {1{`RANDOM}};
  _T_2776_re = _RAND_5172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5173 = {1{`RANDOM}};
  _T_2776_im = _RAND_5173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5174 = {1{`RANDOM}};
  _T_2777_re = _RAND_5174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5175 = {1{`RANDOM}};
  _T_2777_im = _RAND_5175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5176 = {1{`RANDOM}};
  _T_2778_re = _RAND_5176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5177 = {1{`RANDOM}};
  _T_2778_im = _RAND_5177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5178 = {1{`RANDOM}};
  _T_2779_re = _RAND_5178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5179 = {1{`RANDOM}};
  _T_2779_im = _RAND_5179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5180 = {1{`RANDOM}};
  _T_2780_re = _RAND_5180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5181 = {1{`RANDOM}};
  _T_2780_im = _RAND_5181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5182 = {1{`RANDOM}};
  _T_2781_re = _RAND_5182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5183 = {1{`RANDOM}};
  _T_2781_im = _RAND_5183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5184 = {1{`RANDOM}};
  _T_2782_re = _RAND_5184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5185 = {1{`RANDOM}};
  _T_2782_im = _RAND_5185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5186 = {1{`RANDOM}};
  _T_2783_re = _RAND_5186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5187 = {1{`RANDOM}};
  _T_2783_im = _RAND_5187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5188 = {1{`RANDOM}};
  _T_2784_re = _RAND_5188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5189 = {1{`RANDOM}};
  _T_2784_im = _RAND_5189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5190 = {1{`RANDOM}};
  _T_2785_re = _RAND_5190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5191 = {1{`RANDOM}};
  _T_2785_im = _RAND_5191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5192 = {1{`RANDOM}};
  _T_2786_re = _RAND_5192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5193 = {1{`RANDOM}};
  _T_2786_im = _RAND_5193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5194 = {1{`RANDOM}};
  _T_2787_re = _RAND_5194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5195 = {1{`RANDOM}};
  _T_2787_im = _RAND_5195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5196 = {1{`RANDOM}};
  _T_2788_re = _RAND_5196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5197 = {1{`RANDOM}};
  _T_2788_im = _RAND_5197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5198 = {1{`RANDOM}};
  _T_2789_re = _RAND_5198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5199 = {1{`RANDOM}};
  _T_2789_im = _RAND_5199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5200 = {1{`RANDOM}};
  _T_2790_re = _RAND_5200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5201 = {1{`RANDOM}};
  _T_2790_im = _RAND_5201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5202 = {1{`RANDOM}};
  _T_2791_re = _RAND_5202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5203 = {1{`RANDOM}};
  _T_2791_im = _RAND_5203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5204 = {1{`RANDOM}};
  _T_2792_re = _RAND_5204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5205 = {1{`RANDOM}};
  _T_2792_im = _RAND_5205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5206 = {1{`RANDOM}};
  _T_2793_re = _RAND_5206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5207 = {1{`RANDOM}};
  _T_2793_im = _RAND_5207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5208 = {1{`RANDOM}};
  _T_2794_re = _RAND_5208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5209 = {1{`RANDOM}};
  _T_2794_im = _RAND_5209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5210 = {1{`RANDOM}};
  _T_2795_re = _RAND_5210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5211 = {1{`RANDOM}};
  _T_2795_im = _RAND_5211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5212 = {1{`RANDOM}};
  _T_2796_re = _RAND_5212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5213 = {1{`RANDOM}};
  _T_2796_im = _RAND_5213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5214 = {1{`RANDOM}};
  _T_2797_re = _RAND_5214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5215 = {1{`RANDOM}};
  _T_2797_im = _RAND_5215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5216 = {1{`RANDOM}};
  _T_2798_re = _RAND_5216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5217 = {1{`RANDOM}};
  _T_2798_im = _RAND_5217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5218 = {1{`RANDOM}};
  _T_2799_re = _RAND_5218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5219 = {1{`RANDOM}};
  _T_2799_im = _RAND_5219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5220 = {1{`RANDOM}};
  _T_2800_re = _RAND_5220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5221 = {1{`RANDOM}};
  _T_2800_im = _RAND_5221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5222 = {1{`RANDOM}};
  _T_2801_re = _RAND_5222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5223 = {1{`RANDOM}};
  _T_2801_im = _RAND_5223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5224 = {1{`RANDOM}};
  _T_2802_re = _RAND_5224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5225 = {1{`RANDOM}};
  _T_2802_im = _RAND_5225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5226 = {1{`RANDOM}};
  _T_2803_re = _RAND_5226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5227 = {1{`RANDOM}};
  _T_2803_im = _RAND_5227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5228 = {1{`RANDOM}};
  _T_2804_re = _RAND_5228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5229 = {1{`RANDOM}};
  _T_2804_im = _RAND_5229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5230 = {1{`RANDOM}};
  _T_2805_re = _RAND_5230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5231 = {1{`RANDOM}};
  _T_2805_im = _RAND_5231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5232 = {1{`RANDOM}};
  _T_2806_re = _RAND_5232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5233 = {1{`RANDOM}};
  _T_2806_im = _RAND_5233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5234 = {1{`RANDOM}};
  _T_2807_re = _RAND_5234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5235 = {1{`RANDOM}};
  _T_2807_im = _RAND_5235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5236 = {1{`RANDOM}};
  _T_2808_re = _RAND_5236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5237 = {1{`RANDOM}};
  _T_2808_im = _RAND_5237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5238 = {1{`RANDOM}};
  _T_2809_re = _RAND_5238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5239 = {1{`RANDOM}};
  _T_2809_im = _RAND_5239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5240 = {1{`RANDOM}};
  _T_2810_re = _RAND_5240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5241 = {1{`RANDOM}};
  _T_2810_im = _RAND_5241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5242 = {1{`RANDOM}};
  _T_2811_re = _RAND_5242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5243 = {1{`RANDOM}};
  _T_2811_im = _RAND_5243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5244 = {1{`RANDOM}};
  _T_2812_re = _RAND_5244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5245 = {1{`RANDOM}};
  _T_2812_im = _RAND_5245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5246 = {1{`RANDOM}};
  _T_2813_re = _RAND_5246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5247 = {1{`RANDOM}};
  _T_2813_im = _RAND_5247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5248 = {1{`RANDOM}};
  _T_2814_re = _RAND_5248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5249 = {1{`RANDOM}};
  _T_2814_im = _RAND_5249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5250 = {1{`RANDOM}};
  _T_2815_re = _RAND_5250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5251 = {1{`RANDOM}};
  _T_2815_im = _RAND_5251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5252 = {1{`RANDOM}};
  _T_2816_re = _RAND_5252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5253 = {1{`RANDOM}};
  _T_2816_im = _RAND_5253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5254 = {1{`RANDOM}};
  _T_2817_re = _RAND_5254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5255 = {1{`RANDOM}};
  _T_2817_im = _RAND_5255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5256 = {1{`RANDOM}};
  _T_2818_re = _RAND_5256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5257 = {1{`RANDOM}};
  _T_2818_im = _RAND_5257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5258 = {1{`RANDOM}};
  _T_2819_re = _RAND_5258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5259 = {1{`RANDOM}};
  _T_2819_im = _RAND_5259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5260 = {1{`RANDOM}};
  _T_2820_re = _RAND_5260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5261 = {1{`RANDOM}};
  _T_2820_im = _RAND_5261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5262 = {1{`RANDOM}};
  _T_2821_re = _RAND_5262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5263 = {1{`RANDOM}};
  _T_2821_im = _RAND_5263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5264 = {1{`RANDOM}};
  _T_2822_re = _RAND_5264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5265 = {1{`RANDOM}};
  _T_2822_im = _RAND_5265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5266 = {1{`RANDOM}};
  _T_2823_re = _RAND_5266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5267 = {1{`RANDOM}};
  _T_2823_im = _RAND_5267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5268 = {1{`RANDOM}};
  _T_2824_re = _RAND_5268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5269 = {1{`RANDOM}};
  _T_2824_im = _RAND_5269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5270 = {1{`RANDOM}};
  _T_2825_re = _RAND_5270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5271 = {1{`RANDOM}};
  _T_2825_im = _RAND_5271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5272 = {1{`RANDOM}};
  _T_2826_re = _RAND_5272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5273 = {1{`RANDOM}};
  _T_2826_im = _RAND_5273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5274 = {1{`RANDOM}};
  _T_2827_re = _RAND_5274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5275 = {1{`RANDOM}};
  _T_2827_im = _RAND_5275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5276 = {1{`RANDOM}};
  _T_2828_re = _RAND_5276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5277 = {1{`RANDOM}};
  _T_2828_im = _RAND_5277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5278 = {1{`RANDOM}};
  _T_2829_re = _RAND_5278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5279 = {1{`RANDOM}};
  _T_2829_im = _RAND_5279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5280 = {1{`RANDOM}};
  _T_2830_re = _RAND_5280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5281 = {1{`RANDOM}};
  _T_2830_im = _RAND_5281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5282 = {1{`RANDOM}};
  _T_2831_re = _RAND_5282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5283 = {1{`RANDOM}};
  _T_2831_im = _RAND_5283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5284 = {1{`RANDOM}};
  _T_2832_re = _RAND_5284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5285 = {1{`RANDOM}};
  _T_2832_im = _RAND_5285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5286 = {1{`RANDOM}};
  _T_2833_re = _RAND_5286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5287 = {1{`RANDOM}};
  _T_2833_im = _RAND_5287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5288 = {1{`RANDOM}};
  _T_2834_re = _RAND_5288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5289 = {1{`RANDOM}};
  _T_2834_im = _RAND_5289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5290 = {1{`RANDOM}};
  _T_2835_re = _RAND_5290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5291 = {1{`RANDOM}};
  _T_2835_im = _RAND_5291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5292 = {1{`RANDOM}};
  _T_2836_re = _RAND_5292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5293 = {1{`RANDOM}};
  _T_2836_im = _RAND_5293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5294 = {1{`RANDOM}};
  _T_2837_re = _RAND_5294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5295 = {1{`RANDOM}};
  _T_2837_im = _RAND_5295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5296 = {1{`RANDOM}};
  _T_2838_re = _RAND_5296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5297 = {1{`RANDOM}};
  _T_2838_im = _RAND_5297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5298 = {1{`RANDOM}};
  _T_2839_re = _RAND_5298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5299 = {1{`RANDOM}};
  _T_2839_im = _RAND_5299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5300 = {1{`RANDOM}};
  _T_2840_re = _RAND_5300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5301 = {1{`RANDOM}};
  _T_2840_im = _RAND_5301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5302 = {1{`RANDOM}};
  _T_2841_re = _RAND_5302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5303 = {1{`RANDOM}};
  _T_2841_im = _RAND_5303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5304 = {1{`RANDOM}};
  _T_2842_re = _RAND_5304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5305 = {1{`RANDOM}};
  _T_2842_im = _RAND_5305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5306 = {1{`RANDOM}};
  _T_2843_re = _RAND_5306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5307 = {1{`RANDOM}};
  _T_2843_im = _RAND_5307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5308 = {1{`RANDOM}};
  _T_2844_re = _RAND_5308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5309 = {1{`RANDOM}};
  _T_2844_im = _RAND_5309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5310 = {1{`RANDOM}};
  _T_2845_re = _RAND_5310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5311 = {1{`RANDOM}};
  _T_2845_im = _RAND_5311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5312 = {1{`RANDOM}};
  _T_2846_re = _RAND_5312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5313 = {1{`RANDOM}};
  _T_2846_im = _RAND_5313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5314 = {1{`RANDOM}};
  _T_2847_re = _RAND_5314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5315 = {1{`RANDOM}};
  _T_2847_im = _RAND_5315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5316 = {1{`RANDOM}};
  _T_2848_re = _RAND_5316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5317 = {1{`RANDOM}};
  _T_2848_im = _RAND_5317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5318 = {1{`RANDOM}};
  _T_2849_re = _RAND_5318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5319 = {1{`RANDOM}};
  _T_2849_im = _RAND_5319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5320 = {1{`RANDOM}};
  _T_2850_re = _RAND_5320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5321 = {1{`RANDOM}};
  _T_2850_im = _RAND_5321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5322 = {1{`RANDOM}};
  _T_2851_re = _RAND_5322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5323 = {1{`RANDOM}};
  _T_2851_im = _RAND_5323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5324 = {1{`RANDOM}};
  _T_2852_re = _RAND_5324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5325 = {1{`RANDOM}};
  _T_2852_im = _RAND_5325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5326 = {1{`RANDOM}};
  _T_2853_re = _RAND_5326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5327 = {1{`RANDOM}};
  _T_2853_im = _RAND_5327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5328 = {1{`RANDOM}};
  _T_2854_re = _RAND_5328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5329 = {1{`RANDOM}};
  _T_2854_im = _RAND_5329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5330 = {1{`RANDOM}};
  _T_2855_re = _RAND_5330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5331 = {1{`RANDOM}};
  _T_2855_im = _RAND_5331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5332 = {1{`RANDOM}};
  _T_2856_re = _RAND_5332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5333 = {1{`RANDOM}};
  _T_2856_im = _RAND_5333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5334 = {1{`RANDOM}};
  _T_2857_re = _RAND_5334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5335 = {1{`RANDOM}};
  _T_2857_im = _RAND_5335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5336 = {1{`RANDOM}};
  _T_2858_re = _RAND_5336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5337 = {1{`RANDOM}};
  _T_2858_im = _RAND_5337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5338 = {1{`RANDOM}};
  _T_2859_re = _RAND_5338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5339 = {1{`RANDOM}};
  _T_2859_im = _RAND_5339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5340 = {1{`RANDOM}};
  _T_2860_re = _RAND_5340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5341 = {1{`RANDOM}};
  _T_2860_im = _RAND_5341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5342 = {1{`RANDOM}};
  _T_2861_re = _RAND_5342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5343 = {1{`RANDOM}};
  _T_2861_im = _RAND_5343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5344 = {1{`RANDOM}};
  _T_2862_re = _RAND_5344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5345 = {1{`RANDOM}};
  _T_2862_im = _RAND_5345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5346 = {1{`RANDOM}};
  _T_2863_re = _RAND_5346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5347 = {1{`RANDOM}};
  _T_2863_im = _RAND_5347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5348 = {1{`RANDOM}};
  _T_2864_re = _RAND_5348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5349 = {1{`RANDOM}};
  _T_2864_im = _RAND_5349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5350 = {1{`RANDOM}};
  _T_2865_re = _RAND_5350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5351 = {1{`RANDOM}};
  _T_2865_im = _RAND_5351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5352 = {1{`RANDOM}};
  _T_2866_re = _RAND_5352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5353 = {1{`RANDOM}};
  _T_2866_im = _RAND_5353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5354 = {1{`RANDOM}};
  _T_2867_re = _RAND_5354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5355 = {1{`RANDOM}};
  _T_2867_im = _RAND_5355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5356 = {1{`RANDOM}};
  _T_2868_re = _RAND_5356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5357 = {1{`RANDOM}};
  _T_2868_im = _RAND_5357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5358 = {1{`RANDOM}};
  _T_2869_re = _RAND_5358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5359 = {1{`RANDOM}};
  _T_2869_im = _RAND_5359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5360 = {1{`RANDOM}};
  _T_2870_re = _RAND_5360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5361 = {1{`RANDOM}};
  _T_2870_im = _RAND_5361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5362 = {1{`RANDOM}};
  _T_2871_re = _RAND_5362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5363 = {1{`RANDOM}};
  _T_2871_im = _RAND_5363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5364 = {1{`RANDOM}};
  _T_2872_re = _RAND_5364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5365 = {1{`RANDOM}};
  _T_2872_im = _RAND_5365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5366 = {1{`RANDOM}};
  _T_2873_re = _RAND_5366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5367 = {1{`RANDOM}};
  _T_2873_im = _RAND_5367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5368 = {1{`RANDOM}};
  _T_2874_re = _RAND_5368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5369 = {1{`RANDOM}};
  _T_2874_im = _RAND_5369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5370 = {1{`RANDOM}};
  _T_2875_re = _RAND_5370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5371 = {1{`RANDOM}};
  _T_2875_im = _RAND_5371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5372 = {1{`RANDOM}};
  _T_2876_re = _RAND_5372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5373 = {1{`RANDOM}};
  _T_2876_im = _RAND_5373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5374 = {1{`RANDOM}};
  _T_2877_re = _RAND_5374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5375 = {1{`RANDOM}};
  _T_2877_im = _RAND_5375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5376 = {1{`RANDOM}};
  _T_2878_re = _RAND_5376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5377 = {1{`RANDOM}};
  _T_2878_im = _RAND_5377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5378 = {1{`RANDOM}};
  _T_2879_re = _RAND_5378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5379 = {1{`RANDOM}};
  _T_2879_im = _RAND_5379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5380 = {1{`RANDOM}};
  _T_2880_re = _RAND_5380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5381 = {1{`RANDOM}};
  _T_2880_im = _RAND_5381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5382 = {1{`RANDOM}};
  _T_2881_re = _RAND_5382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5383 = {1{`RANDOM}};
  _T_2881_im = _RAND_5383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5384 = {1{`RANDOM}};
  _T_2882_re = _RAND_5384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5385 = {1{`RANDOM}};
  _T_2882_im = _RAND_5385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5386 = {1{`RANDOM}};
  _T_2883_re = _RAND_5386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5387 = {1{`RANDOM}};
  _T_2883_im = _RAND_5387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5388 = {1{`RANDOM}};
  _T_2884_re = _RAND_5388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5389 = {1{`RANDOM}};
  _T_2884_im = _RAND_5389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5390 = {1{`RANDOM}};
  _T_2885_re = _RAND_5390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5391 = {1{`RANDOM}};
  _T_2885_im = _RAND_5391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5392 = {1{`RANDOM}};
  _T_2886_re = _RAND_5392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5393 = {1{`RANDOM}};
  _T_2886_im = _RAND_5393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5394 = {1{`RANDOM}};
  _T_2887_re = _RAND_5394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5395 = {1{`RANDOM}};
  _T_2887_im = _RAND_5395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5396 = {1{`RANDOM}};
  _T_2888_re = _RAND_5396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5397 = {1{`RANDOM}};
  _T_2888_im = _RAND_5397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5398 = {1{`RANDOM}};
  _T_2889_re = _RAND_5398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5399 = {1{`RANDOM}};
  _T_2889_im = _RAND_5399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5400 = {1{`RANDOM}};
  _T_2890_re = _RAND_5400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5401 = {1{`RANDOM}};
  _T_2890_im = _RAND_5401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5402 = {1{`RANDOM}};
  _T_2891_re = _RAND_5402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5403 = {1{`RANDOM}};
  _T_2891_im = _RAND_5403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5404 = {1{`RANDOM}};
  _T_2892_re = _RAND_5404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5405 = {1{`RANDOM}};
  _T_2892_im = _RAND_5405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5406 = {1{`RANDOM}};
  _T_2893_re = _RAND_5406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5407 = {1{`RANDOM}};
  _T_2893_im = _RAND_5407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5408 = {1{`RANDOM}};
  _T_2894_re = _RAND_5408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5409 = {1{`RANDOM}};
  _T_2894_im = _RAND_5409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5410 = {1{`RANDOM}};
  _T_2895_re = _RAND_5410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5411 = {1{`RANDOM}};
  _T_2895_im = _RAND_5411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5412 = {1{`RANDOM}};
  _T_2896_re = _RAND_5412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5413 = {1{`RANDOM}};
  _T_2896_im = _RAND_5413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5414 = {1{`RANDOM}};
  _T_2897_re = _RAND_5414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5415 = {1{`RANDOM}};
  _T_2897_im = _RAND_5415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5416 = {1{`RANDOM}};
  _T_2898_re = _RAND_5416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5417 = {1{`RANDOM}};
  _T_2898_im = _RAND_5417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5418 = {1{`RANDOM}};
  _T_2899_re = _RAND_5418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5419 = {1{`RANDOM}};
  _T_2899_im = _RAND_5419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5420 = {1{`RANDOM}};
  _T_2900_re = _RAND_5420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5421 = {1{`RANDOM}};
  _T_2900_im = _RAND_5421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5422 = {1{`RANDOM}};
  _T_2901_re = _RAND_5422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5423 = {1{`RANDOM}};
  _T_2901_im = _RAND_5423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5424 = {1{`RANDOM}};
  _T_2902_re = _RAND_5424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5425 = {1{`RANDOM}};
  _T_2902_im = _RAND_5425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5426 = {1{`RANDOM}};
  _T_2903_re = _RAND_5426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5427 = {1{`RANDOM}};
  _T_2903_im = _RAND_5427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5428 = {1{`RANDOM}};
  _T_2904_re = _RAND_5428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5429 = {1{`RANDOM}};
  _T_2904_im = _RAND_5429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5430 = {1{`RANDOM}};
  _T_2905_re = _RAND_5430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5431 = {1{`RANDOM}};
  _T_2905_im = _RAND_5431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5432 = {1{`RANDOM}};
  _T_2906_re = _RAND_5432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5433 = {1{`RANDOM}};
  _T_2906_im = _RAND_5433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5434 = {1{`RANDOM}};
  _T_2907_re = _RAND_5434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5435 = {1{`RANDOM}};
  _T_2907_im = _RAND_5435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5436 = {1{`RANDOM}};
  _T_2908_re = _RAND_5436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5437 = {1{`RANDOM}};
  _T_2908_im = _RAND_5437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5438 = {1{`RANDOM}};
  _T_2909_re = _RAND_5438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5439 = {1{`RANDOM}};
  _T_2909_im = _RAND_5439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5440 = {1{`RANDOM}};
  _T_2910_re = _RAND_5440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5441 = {1{`RANDOM}};
  _T_2910_im = _RAND_5441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5442 = {1{`RANDOM}};
  _T_2911_re = _RAND_5442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5443 = {1{`RANDOM}};
  _T_2911_im = _RAND_5443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5444 = {1{`RANDOM}};
  _T_2912_re = _RAND_5444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5445 = {1{`RANDOM}};
  _T_2912_im = _RAND_5445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5446 = {1{`RANDOM}};
  _T_2913_re = _RAND_5446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5447 = {1{`RANDOM}};
  _T_2913_im = _RAND_5447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5448 = {1{`RANDOM}};
  _T_2914_re = _RAND_5448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5449 = {1{`RANDOM}};
  _T_2914_im = _RAND_5449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5450 = {1{`RANDOM}};
  _T_2915_re = _RAND_5450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5451 = {1{`RANDOM}};
  _T_2915_im = _RAND_5451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5452 = {1{`RANDOM}};
  _T_2916_re = _RAND_5452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5453 = {1{`RANDOM}};
  _T_2916_im = _RAND_5453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5454 = {1{`RANDOM}};
  _T_2917_re = _RAND_5454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5455 = {1{`RANDOM}};
  _T_2917_im = _RAND_5455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5456 = {1{`RANDOM}};
  _T_2918_re = _RAND_5456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5457 = {1{`RANDOM}};
  _T_2918_im = _RAND_5457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5458 = {1{`RANDOM}};
  _T_2919_re = _RAND_5458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5459 = {1{`RANDOM}};
  _T_2919_im = _RAND_5459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5460 = {1{`RANDOM}};
  _T_2920_re = _RAND_5460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5461 = {1{`RANDOM}};
  _T_2920_im = _RAND_5461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5462 = {1{`RANDOM}};
  _T_2921_re = _RAND_5462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5463 = {1{`RANDOM}};
  _T_2921_im = _RAND_5463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5464 = {1{`RANDOM}};
  _T_2922_re = _RAND_5464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5465 = {1{`RANDOM}};
  _T_2922_im = _RAND_5465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5466 = {1{`RANDOM}};
  _T_2923_re = _RAND_5466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5467 = {1{`RANDOM}};
  _T_2923_im = _RAND_5467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5468 = {1{`RANDOM}};
  _T_2924_re = _RAND_5468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5469 = {1{`RANDOM}};
  _T_2924_im = _RAND_5469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5470 = {1{`RANDOM}};
  _T_2925_re = _RAND_5470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5471 = {1{`RANDOM}};
  _T_2925_im = _RAND_5471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5472 = {1{`RANDOM}};
  _T_2926_re = _RAND_5472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5473 = {1{`RANDOM}};
  _T_2926_im = _RAND_5473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5474 = {1{`RANDOM}};
  _T_2927_re = _RAND_5474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5475 = {1{`RANDOM}};
  _T_2927_im = _RAND_5475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5476 = {1{`RANDOM}};
  _T_2928_re = _RAND_5476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5477 = {1{`RANDOM}};
  _T_2928_im = _RAND_5477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5478 = {1{`RANDOM}};
  _T_2929_re = _RAND_5478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5479 = {1{`RANDOM}};
  _T_2929_im = _RAND_5479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5480 = {1{`RANDOM}};
  _T_2930_re = _RAND_5480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5481 = {1{`RANDOM}};
  _T_2930_im = _RAND_5481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5482 = {1{`RANDOM}};
  _T_2931_re = _RAND_5482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5483 = {1{`RANDOM}};
  _T_2931_im = _RAND_5483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5484 = {1{`RANDOM}};
  _T_2932_re = _RAND_5484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5485 = {1{`RANDOM}};
  _T_2932_im = _RAND_5485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5486 = {1{`RANDOM}};
  _T_2933_re = _RAND_5486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5487 = {1{`RANDOM}};
  _T_2933_im = _RAND_5487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5488 = {1{`RANDOM}};
  _T_2934_re = _RAND_5488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5489 = {1{`RANDOM}};
  _T_2934_im = _RAND_5489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5490 = {1{`RANDOM}};
  _T_2935_re = _RAND_5490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5491 = {1{`RANDOM}};
  _T_2935_im = _RAND_5491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5492 = {1{`RANDOM}};
  _T_2936_re = _RAND_5492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5493 = {1{`RANDOM}};
  _T_2936_im = _RAND_5493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5494 = {1{`RANDOM}};
  _T_2937_re = _RAND_5494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5495 = {1{`RANDOM}};
  _T_2937_im = _RAND_5495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5496 = {1{`RANDOM}};
  _T_2938_re = _RAND_5496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5497 = {1{`RANDOM}};
  _T_2938_im = _RAND_5497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5498 = {1{`RANDOM}};
  _T_2939_re = _RAND_5498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5499 = {1{`RANDOM}};
  _T_2939_im = _RAND_5499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5500 = {1{`RANDOM}};
  _T_2940_re = _RAND_5500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5501 = {1{`RANDOM}};
  _T_2940_im = _RAND_5501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5502 = {1{`RANDOM}};
  _T_2941_re = _RAND_5502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5503 = {1{`RANDOM}};
  _T_2941_im = _RAND_5503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5504 = {1{`RANDOM}};
  _T_2942_re = _RAND_5504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5505 = {1{`RANDOM}};
  _T_2942_im = _RAND_5505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5506 = {1{`RANDOM}};
  _T_2943_re = _RAND_5506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5507 = {1{`RANDOM}};
  _T_2943_im = _RAND_5507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5508 = {1{`RANDOM}};
  _T_2944_re = _RAND_5508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5509 = {1{`RANDOM}};
  _T_2944_im = _RAND_5509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5510 = {1{`RANDOM}};
  _T_2945_re = _RAND_5510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5511 = {1{`RANDOM}};
  _T_2945_im = _RAND_5511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5512 = {1{`RANDOM}};
  _T_2946_re = _RAND_5512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5513 = {1{`RANDOM}};
  _T_2946_im = _RAND_5513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5514 = {1{`RANDOM}};
  _T_2947_re = _RAND_5514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5515 = {1{`RANDOM}};
  _T_2947_im = _RAND_5515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5516 = {1{`RANDOM}};
  _T_2948_re = _RAND_5516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5517 = {1{`RANDOM}};
  _T_2948_im = _RAND_5517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5518 = {1{`RANDOM}};
  _T_2949_re = _RAND_5518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5519 = {1{`RANDOM}};
  _T_2949_im = _RAND_5519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5520 = {1{`RANDOM}};
  _T_2950_re = _RAND_5520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5521 = {1{`RANDOM}};
  _T_2950_im = _RAND_5521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5522 = {1{`RANDOM}};
  _T_2951_re = _RAND_5522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5523 = {1{`RANDOM}};
  _T_2951_im = _RAND_5523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5524 = {1{`RANDOM}};
  _T_2952_re = _RAND_5524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5525 = {1{`RANDOM}};
  _T_2952_im = _RAND_5525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5526 = {1{`RANDOM}};
  _T_2953_re = _RAND_5526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5527 = {1{`RANDOM}};
  _T_2953_im = _RAND_5527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5528 = {1{`RANDOM}};
  _T_2954_re = _RAND_5528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5529 = {1{`RANDOM}};
  _T_2954_im = _RAND_5529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5530 = {1{`RANDOM}};
  _T_2955_re = _RAND_5530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5531 = {1{`RANDOM}};
  _T_2955_im = _RAND_5531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5532 = {1{`RANDOM}};
  _T_2956_re = _RAND_5532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5533 = {1{`RANDOM}};
  _T_2956_im = _RAND_5533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5534 = {1{`RANDOM}};
  _T_2957_re = _RAND_5534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5535 = {1{`RANDOM}};
  _T_2957_im = _RAND_5535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5536 = {1{`RANDOM}};
  _T_2958_re = _RAND_5536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5537 = {1{`RANDOM}};
  _T_2958_im = _RAND_5537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5538 = {1{`RANDOM}};
  _T_2959_re = _RAND_5538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5539 = {1{`RANDOM}};
  _T_2959_im = _RAND_5539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5540 = {1{`RANDOM}};
  _T_2960_re = _RAND_5540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5541 = {1{`RANDOM}};
  _T_2960_im = _RAND_5541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5542 = {1{`RANDOM}};
  _T_2961_re = _RAND_5542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5543 = {1{`RANDOM}};
  _T_2961_im = _RAND_5543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5544 = {1{`RANDOM}};
  _T_2962_re = _RAND_5544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5545 = {1{`RANDOM}};
  _T_2962_im = _RAND_5545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5546 = {1{`RANDOM}};
  _T_2963_re = _RAND_5546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5547 = {1{`RANDOM}};
  _T_2963_im = _RAND_5547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5548 = {1{`RANDOM}};
  _T_2964_re = _RAND_5548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5549 = {1{`RANDOM}};
  _T_2964_im = _RAND_5549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5550 = {1{`RANDOM}};
  _T_2965_re = _RAND_5550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5551 = {1{`RANDOM}};
  _T_2965_im = _RAND_5551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5552 = {1{`RANDOM}};
  _T_2966_re = _RAND_5552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5553 = {1{`RANDOM}};
  _T_2966_im = _RAND_5553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5554 = {1{`RANDOM}};
  _T_2967_re = _RAND_5554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5555 = {1{`RANDOM}};
  _T_2967_im = _RAND_5555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5556 = {1{`RANDOM}};
  _T_2968_re = _RAND_5556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5557 = {1{`RANDOM}};
  _T_2968_im = _RAND_5557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5558 = {1{`RANDOM}};
  _T_2969_re = _RAND_5558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5559 = {1{`RANDOM}};
  _T_2969_im = _RAND_5559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5560 = {1{`RANDOM}};
  _T_2970_re = _RAND_5560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5561 = {1{`RANDOM}};
  _T_2970_im = _RAND_5561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5562 = {1{`RANDOM}};
  _T_2971_re = _RAND_5562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5563 = {1{`RANDOM}};
  _T_2971_im = _RAND_5563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5564 = {1{`RANDOM}};
  _T_2972_re = _RAND_5564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5565 = {1{`RANDOM}};
  _T_2972_im = _RAND_5565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5566 = {1{`RANDOM}};
  _T_2973_re = _RAND_5566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5567 = {1{`RANDOM}};
  _T_2973_im = _RAND_5567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5568 = {1{`RANDOM}};
  _T_2974_re = _RAND_5568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5569 = {1{`RANDOM}};
  _T_2974_im = _RAND_5569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5570 = {1{`RANDOM}};
  _T_2975_re = _RAND_5570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5571 = {1{`RANDOM}};
  _T_2975_im = _RAND_5571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5572 = {1{`RANDOM}};
  _T_2976_re = _RAND_5572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5573 = {1{`RANDOM}};
  _T_2976_im = _RAND_5573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5574 = {1{`RANDOM}};
  _T_2977_re = _RAND_5574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5575 = {1{`RANDOM}};
  _T_2977_im = _RAND_5575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5576 = {1{`RANDOM}};
  _T_2978_re = _RAND_5576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5577 = {1{`RANDOM}};
  _T_2978_im = _RAND_5577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5578 = {1{`RANDOM}};
  _T_2979_re = _RAND_5578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5579 = {1{`RANDOM}};
  _T_2979_im = _RAND_5579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5580 = {1{`RANDOM}};
  _T_2980_re = _RAND_5580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5581 = {1{`RANDOM}};
  _T_2980_im = _RAND_5581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5582 = {1{`RANDOM}};
  _T_2981_re = _RAND_5582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5583 = {1{`RANDOM}};
  _T_2981_im = _RAND_5583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5584 = {1{`RANDOM}};
  _T_2982_re = _RAND_5584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5585 = {1{`RANDOM}};
  _T_2982_im = _RAND_5585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5586 = {1{`RANDOM}};
  _T_2983_re = _RAND_5586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5587 = {1{`RANDOM}};
  _T_2983_im = _RAND_5587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5588 = {1{`RANDOM}};
  _T_2984_re = _RAND_5588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5589 = {1{`RANDOM}};
  _T_2984_im = _RAND_5589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5590 = {1{`RANDOM}};
  _T_2985_re = _RAND_5590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5591 = {1{`RANDOM}};
  _T_2985_im = _RAND_5591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5592 = {1{`RANDOM}};
  _T_2986_re = _RAND_5592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5593 = {1{`RANDOM}};
  _T_2986_im = _RAND_5593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5594 = {1{`RANDOM}};
  _T_2987_re = _RAND_5594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5595 = {1{`RANDOM}};
  _T_2987_im = _RAND_5595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5596 = {1{`RANDOM}};
  _T_2988_re = _RAND_5596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5597 = {1{`RANDOM}};
  _T_2988_im = _RAND_5597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5598 = {1{`RANDOM}};
  _T_2989_re = _RAND_5598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5599 = {1{`RANDOM}};
  _T_2989_im = _RAND_5599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5600 = {1{`RANDOM}};
  _T_2990_re = _RAND_5600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5601 = {1{`RANDOM}};
  _T_2990_im = _RAND_5601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5602 = {1{`RANDOM}};
  _T_2991_re = _RAND_5602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5603 = {1{`RANDOM}};
  _T_2991_im = _RAND_5603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5604 = {1{`RANDOM}};
  _T_2992_re = _RAND_5604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5605 = {1{`RANDOM}};
  _T_2992_im = _RAND_5605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5606 = {1{`RANDOM}};
  _T_2993_re = _RAND_5606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5607 = {1{`RANDOM}};
  _T_2993_im = _RAND_5607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5608 = {1{`RANDOM}};
  _T_2994_re = _RAND_5608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5609 = {1{`RANDOM}};
  _T_2994_im = _RAND_5609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5610 = {1{`RANDOM}};
  _T_2995_re = _RAND_5610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5611 = {1{`RANDOM}};
  _T_2995_im = _RAND_5611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5612 = {1{`RANDOM}};
  _T_2996_re = _RAND_5612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5613 = {1{`RANDOM}};
  _T_2996_im = _RAND_5613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5614 = {1{`RANDOM}};
  _T_2997_re = _RAND_5614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5615 = {1{`RANDOM}};
  _T_2997_im = _RAND_5615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5616 = {1{`RANDOM}};
  _T_2998_re = _RAND_5616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5617 = {1{`RANDOM}};
  _T_2998_im = _RAND_5617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5618 = {1{`RANDOM}};
  _T_2999_re = _RAND_5618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5619 = {1{`RANDOM}};
  _T_2999_im = _RAND_5619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5620 = {1{`RANDOM}};
  _T_3000_re = _RAND_5620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5621 = {1{`RANDOM}};
  _T_3000_im = _RAND_5621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5622 = {1{`RANDOM}};
  _T_3001_re = _RAND_5622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5623 = {1{`RANDOM}};
  _T_3001_im = _RAND_5623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5624 = {1{`RANDOM}};
  _T_3002_re = _RAND_5624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5625 = {1{`RANDOM}};
  _T_3002_im = _RAND_5625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5626 = {1{`RANDOM}};
  _T_3003_re = _RAND_5626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5627 = {1{`RANDOM}};
  _T_3003_im = _RAND_5627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5628 = {1{`RANDOM}};
  _T_3004_re = _RAND_5628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5629 = {1{`RANDOM}};
  _T_3004_im = _RAND_5629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5630 = {1{`RANDOM}};
  _T_3005_re = _RAND_5630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5631 = {1{`RANDOM}};
  _T_3005_im = _RAND_5631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5632 = {1{`RANDOM}};
  _T_3006_re = _RAND_5632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5633 = {1{`RANDOM}};
  _T_3006_im = _RAND_5633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5634 = {1{`RANDOM}};
  _T_3007_re = _RAND_5634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5635 = {1{`RANDOM}};
  _T_3007_im = _RAND_5635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5636 = {1{`RANDOM}};
  _T_3008_re = _RAND_5636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5637 = {1{`RANDOM}};
  _T_3008_im = _RAND_5637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5638 = {1{`RANDOM}};
  _T_3009_re = _RAND_5638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5639 = {1{`RANDOM}};
  _T_3009_im = _RAND_5639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5640 = {1{`RANDOM}};
  _T_3010_re = _RAND_5640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5641 = {1{`RANDOM}};
  _T_3010_im = _RAND_5641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5642 = {1{`RANDOM}};
  _T_3011_re = _RAND_5642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5643 = {1{`RANDOM}};
  _T_3011_im = _RAND_5643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5644 = {1{`RANDOM}};
  _T_3012_re = _RAND_5644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5645 = {1{`RANDOM}};
  _T_3012_im = _RAND_5645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5646 = {1{`RANDOM}};
  _T_3013_re = _RAND_5646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5647 = {1{`RANDOM}};
  _T_3013_im = _RAND_5647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5648 = {1{`RANDOM}};
  _T_3014_re = _RAND_5648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5649 = {1{`RANDOM}};
  _T_3014_im = _RAND_5649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5650 = {1{`RANDOM}};
  _T_3015_re = _RAND_5650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5651 = {1{`RANDOM}};
  _T_3015_im = _RAND_5651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5652 = {1{`RANDOM}};
  _T_3016_re = _RAND_5652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5653 = {1{`RANDOM}};
  _T_3016_im = _RAND_5653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5654 = {1{`RANDOM}};
  _T_3017_re = _RAND_5654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5655 = {1{`RANDOM}};
  _T_3017_im = _RAND_5655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5656 = {1{`RANDOM}};
  _T_3018_re = _RAND_5656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5657 = {1{`RANDOM}};
  _T_3018_im = _RAND_5657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5658 = {1{`RANDOM}};
  _T_3019_re = _RAND_5658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5659 = {1{`RANDOM}};
  _T_3019_im = _RAND_5659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5660 = {1{`RANDOM}};
  _T_3020_re = _RAND_5660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5661 = {1{`RANDOM}};
  _T_3020_im = _RAND_5661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5662 = {1{`RANDOM}};
  _T_3021_re = _RAND_5662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5663 = {1{`RANDOM}};
  _T_3021_im = _RAND_5663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5664 = {1{`RANDOM}};
  _T_3022_re = _RAND_5664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5665 = {1{`RANDOM}};
  _T_3022_im = _RAND_5665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5666 = {1{`RANDOM}};
  _T_3023_re = _RAND_5666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5667 = {1{`RANDOM}};
  _T_3023_im = _RAND_5667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5668 = {1{`RANDOM}};
  _T_3024_re = _RAND_5668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5669 = {1{`RANDOM}};
  _T_3024_im = _RAND_5669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5670 = {1{`RANDOM}};
  _T_3025_re = _RAND_5670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5671 = {1{`RANDOM}};
  _T_3025_im = _RAND_5671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5672 = {1{`RANDOM}};
  _T_3026_re = _RAND_5672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5673 = {1{`RANDOM}};
  _T_3026_im = _RAND_5673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5674 = {1{`RANDOM}};
  _T_3027_re = _RAND_5674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5675 = {1{`RANDOM}};
  _T_3027_im = _RAND_5675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5676 = {1{`RANDOM}};
  _T_3028_re = _RAND_5676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5677 = {1{`RANDOM}};
  _T_3028_im = _RAND_5677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5678 = {1{`RANDOM}};
  _T_3029_re = _RAND_5678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5679 = {1{`RANDOM}};
  _T_3029_im = _RAND_5679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5680 = {1{`RANDOM}};
  _T_3030_re = _RAND_5680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5681 = {1{`RANDOM}};
  _T_3030_im = _RAND_5681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5682 = {1{`RANDOM}};
  _T_3031_re = _RAND_5682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5683 = {1{`RANDOM}};
  _T_3031_im = _RAND_5683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5684 = {1{`RANDOM}};
  _T_3032_re = _RAND_5684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5685 = {1{`RANDOM}};
  _T_3032_im = _RAND_5685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5686 = {1{`RANDOM}};
  _T_3033_re = _RAND_5686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5687 = {1{`RANDOM}};
  _T_3033_im = _RAND_5687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5688 = {1{`RANDOM}};
  _T_3034_re = _RAND_5688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5689 = {1{`RANDOM}};
  _T_3034_im = _RAND_5689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5690 = {1{`RANDOM}};
  _T_3035_re = _RAND_5690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5691 = {1{`RANDOM}};
  _T_3035_im = _RAND_5691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5692 = {1{`RANDOM}};
  _T_3036_re = _RAND_5692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5693 = {1{`RANDOM}};
  _T_3036_im = _RAND_5693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5694 = {1{`RANDOM}};
  _T_3037_re = _RAND_5694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5695 = {1{`RANDOM}};
  _T_3037_im = _RAND_5695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5696 = {1{`RANDOM}};
  _T_3038_re = _RAND_5696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5697 = {1{`RANDOM}};
  _T_3038_im = _RAND_5697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5698 = {1{`RANDOM}};
  _T_3039_re = _RAND_5698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5699 = {1{`RANDOM}};
  _T_3039_im = _RAND_5699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5700 = {1{`RANDOM}};
  _T_3040_re = _RAND_5700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5701 = {1{`RANDOM}};
  _T_3040_im = _RAND_5701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5702 = {1{`RANDOM}};
  _T_3041_re = _RAND_5702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5703 = {1{`RANDOM}};
  _T_3041_im = _RAND_5703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5704 = {1{`RANDOM}};
  _T_3042_re = _RAND_5704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5705 = {1{`RANDOM}};
  _T_3042_im = _RAND_5705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5706 = {1{`RANDOM}};
  _T_3043_re = _RAND_5706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5707 = {1{`RANDOM}};
  _T_3043_im = _RAND_5707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5708 = {1{`RANDOM}};
  _T_3044_re = _RAND_5708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5709 = {1{`RANDOM}};
  _T_3044_im = _RAND_5709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5710 = {1{`RANDOM}};
  _T_3045_re = _RAND_5710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5711 = {1{`RANDOM}};
  _T_3045_im = _RAND_5711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5712 = {1{`RANDOM}};
  _T_3046_re = _RAND_5712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5713 = {1{`RANDOM}};
  _T_3046_im = _RAND_5713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5714 = {1{`RANDOM}};
  _T_3047_re = _RAND_5714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5715 = {1{`RANDOM}};
  _T_3047_im = _RAND_5715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5716 = {1{`RANDOM}};
  _T_3048_re = _RAND_5716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5717 = {1{`RANDOM}};
  _T_3048_im = _RAND_5717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5718 = {1{`RANDOM}};
  _T_3049_re = _RAND_5718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5719 = {1{`RANDOM}};
  _T_3049_im = _RAND_5719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5720 = {1{`RANDOM}};
  _T_3050_re = _RAND_5720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5721 = {1{`RANDOM}};
  _T_3050_im = _RAND_5721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5722 = {1{`RANDOM}};
  _T_3051_re = _RAND_5722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5723 = {1{`RANDOM}};
  _T_3051_im = _RAND_5723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5724 = {1{`RANDOM}};
  _T_3052_re = _RAND_5724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5725 = {1{`RANDOM}};
  _T_3052_im = _RAND_5725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5726 = {1{`RANDOM}};
  _T_3053_re = _RAND_5726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5727 = {1{`RANDOM}};
  _T_3053_im = _RAND_5727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5728 = {1{`RANDOM}};
  _T_3054_re = _RAND_5728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5729 = {1{`RANDOM}};
  _T_3054_im = _RAND_5729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5730 = {1{`RANDOM}};
  _T_3055_re = _RAND_5730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5731 = {1{`RANDOM}};
  _T_3055_im = _RAND_5731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5732 = {1{`RANDOM}};
  _T_3056_re = _RAND_5732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5733 = {1{`RANDOM}};
  _T_3056_im = _RAND_5733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5734 = {1{`RANDOM}};
  _T_3057_re = _RAND_5734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5735 = {1{`RANDOM}};
  _T_3057_im = _RAND_5735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5736 = {1{`RANDOM}};
  _T_3058_re = _RAND_5736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5737 = {1{`RANDOM}};
  _T_3058_im = _RAND_5737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5738 = {1{`RANDOM}};
  _T_3059_re = _RAND_5738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5739 = {1{`RANDOM}};
  _T_3059_im = _RAND_5739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5740 = {1{`RANDOM}};
  _T_3060_re = _RAND_5740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5741 = {1{`RANDOM}};
  _T_3060_im = _RAND_5741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5742 = {1{`RANDOM}};
  _T_3061_re = _RAND_5742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5743 = {1{`RANDOM}};
  _T_3061_im = _RAND_5743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5744 = {1{`RANDOM}};
  _T_3062_re = _RAND_5744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5745 = {1{`RANDOM}};
  _T_3062_im = _RAND_5745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5746 = {1{`RANDOM}};
  _T_3063_re = _RAND_5746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5747 = {1{`RANDOM}};
  _T_3063_im = _RAND_5747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5748 = {1{`RANDOM}};
  _T_3064_re = _RAND_5748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5749 = {1{`RANDOM}};
  _T_3064_im = _RAND_5749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5750 = {1{`RANDOM}};
  _T_3065_re = _RAND_5750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5751 = {1{`RANDOM}};
  _T_3065_im = _RAND_5751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5752 = {1{`RANDOM}};
  _T_3066_re = _RAND_5752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5753 = {1{`RANDOM}};
  _T_3066_im = _RAND_5753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5754 = {1{`RANDOM}};
  _T_3067_re = _RAND_5754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5755 = {1{`RANDOM}};
  _T_3067_im = _RAND_5755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5756 = {1{`RANDOM}};
  _T_3068_re = _RAND_5756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5757 = {1{`RANDOM}};
  _T_3068_im = _RAND_5757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5758 = {1{`RANDOM}};
  _T_3069_re = _RAND_5758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5759 = {1{`RANDOM}};
  _T_3069_im = _RAND_5759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5760 = {1{`RANDOM}};
  _T_3070_re = _RAND_5760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5761 = {1{`RANDOM}};
  _T_3070_im = _RAND_5761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5762 = {1{`RANDOM}};
  _T_3071_re = _RAND_5762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5763 = {1{`RANDOM}};
  _T_3071_im = _RAND_5763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5764 = {1{`RANDOM}};
  _T_3072_re = _RAND_5764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5765 = {1{`RANDOM}};
  _T_3072_im = _RAND_5765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5766 = {1{`RANDOM}};
  _T_3073_re = _RAND_5766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5767 = {1{`RANDOM}};
  _T_3073_im = _RAND_5767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5768 = {1{`RANDOM}};
  _T_3074_re = _RAND_5768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5769 = {1{`RANDOM}};
  _T_3074_im = _RAND_5769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5770 = {1{`RANDOM}};
  _T_3075_re = _RAND_5770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5771 = {1{`RANDOM}};
  _T_3075_im = _RAND_5771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5772 = {1{`RANDOM}};
  _T_3076_re = _RAND_5772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5773 = {1{`RANDOM}};
  _T_3076_im = _RAND_5773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5774 = {1{`RANDOM}};
  _T_3077_re = _RAND_5774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5775 = {1{`RANDOM}};
  _T_3077_im = _RAND_5775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5776 = {1{`RANDOM}};
  _T_3078_re = _RAND_5776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5777 = {1{`RANDOM}};
  _T_3078_im = _RAND_5777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5778 = {1{`RANDOM}};
  _T_3079_re = _RAND_5778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5779 = {1{`RANDOM}};
  _T_3079_im = _RAND_5779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5780 = {1{`RANDOM}};
  _T_3080_re = _RAND_5780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5781 = {1{`RANDOM}};
  _T_3080_im = _RAND_5781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5782 = {1{`RANDOM}};
  _T_3081_re = _RAND_5782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5783 = {1{`RANDOM}};
  _T_3081_im = _RAND_5783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5784 = {1{`RANDOM}};
  _T_3082_re = _RAND_5784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5785 = {1{`RANDOM}};
  _T_3082_im = _RAND_5785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5786 = {1{`RANDOM}};
  _T_3083_re = _RAND_5786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5787 = {1{`RANDOM}};
  _T_3083_im = _RAND_5787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5788 = {1{`RANDOM}};
  _T_3084_re = _RAND_5788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5789 = {1{`RANDOM}};
  _T_3084_im = _RAND_5789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5790 = {1{`RANDOM}};
  _T_3085_re = _RAND_5790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5791 = {1{`RANDOM}};
  _T_3085_im = _RAND_5791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5792 = {1{`RANDOM}};
  _T_3086_re = _RAND_5792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5793 = {1{`RANDOM}};
  _T_3086_im = _RAND_5793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5794 = {1{`RANDOM}};
  _T_3087_re = _RAND_5794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5795 = {1{`RANDOM}};
  _T_3087_im = _RAND_5795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5796 = {1{`RANDOM}};
  _T_3088_re = _RAND_5796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5797 = {1{`RANDOM}};
  _T_3088_im = _RAND_5797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5798 = {1{`RANDOM}};
  _T_3089_re = _RAND_5798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5799 = {1{`RANDOM}};
  _T_3089_im = _RAND_5799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5800 = {1{`RANDOM}};
  _T_3090_re = _RAND_5800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5801 = {1{`RANDOM}};
  _T_3090_im = _RAND_5801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5802 = {1{`RANDOM}};
  _T_3091_re = _RAND_5802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5803 = {1{`RANDOM}};
  _T_3091_im = _RAND_5803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5804 = {1{`RANDOM}};
  _T_3092_re = _RAND_5804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5805 = {1{`RANDOM}};
  _T_3092_im = _RAND_5805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5806 = {1{`RANDOM}};
  _T_3093_re = _RAND_5806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5807 = {1{`RANDOM}};
  _T_3093_im = _RAND_5807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5808 = {1{`RANDOM}};
  _T_3094_re = _RAND_5808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5809 = {1{`RANDOM}};
  _T_3094_im = _RAND_5809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5810 = {1{`RANDOM}};
  _T_3095_re = _RAND_5810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5811 = {1{`RANDOM}};
  _T_3095_im = _RAND_5811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5812 = {1{`RANDOM}};
  _T_3096_re = _RAND_5812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5813 = {1{`RANDOM}};
  _T_3096_im = _RAND_5813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5814 = {1{`RANDOM}};
  _T_3097_re = _RAND_5814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5815 = {1{`RANDOM}};
  _T_3097_im = _RAND_5815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5816 = {1{`RANDOM}};
  _T_3098_re = _RAND_5816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5817 = {1{`RANDOM}};
  _T_3098_im = _RAND_5817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5818 = {1{`RANDOM}};
  _T_3099_re = _RAND_5818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5819 = {1{`RANDOM}};
  _T_3099_im = _RAND_5819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5820 = {1{`RANDOM}};
  _T_3100_re = _RAND_5820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5821 = {1{`RANDOM}};
  _T_3100_im = _RAND_5821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5822 = {1{`RANDOM}};
  _T_3101_re = _RAND_5822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5823 = {1{`RANDOM}};
  _T_3101_im = _RAND_5823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5824 = {1{`RANDOM}};
  _T_3102_re = _RAND_5824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5825 = {1{`RANDOM}};
  _T_3102_im = _RAND_5825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5826 = {1{`RANDOM}};
  _T_3103_re = _RAND_5826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5827 = {1{`RANDOM}};
  _T_3103_im = _RAND_5827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5828 = {1{`RANDOM}};
  _T_3104_re = _RAND_5828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5829 = {1{`RANDOM}};
  _T_3104_im = _RAND_5829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5830 = {1{`RANDOM}};
  _T_3105_re = _RAND_5830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5831 = {1{`RANDOM}};
  _T_3105_im = _RAND_5831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5832 = {1{`RANDOM}};
  _T_3106_re = _RAND_5832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5833 = {1{`RANDOM}};
  _T_3106_im = _RAND_5833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5834 = {1{`RANDOM}};
  _T_3107_re = _RAND_5834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5835 = {1{`RANDOM}};
  _T_3107_im = _RAND_5835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5836 = {1{`RANDOM}};
  _T_3108_re = _RAND_5836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5837 = {1{`RANDOM}};
  _T_3108_im = _RAND_5837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5838 = {1{`RANDOM}};
  _T_3109_re = _RAND_5838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5839 = {1{`RANDOM}};
  _T_3109_im = _RAND_5839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5840 = {1{`RANDOM}};
  _T_3110_re = _RAND_5840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5841 = {1{`RANDOM}};
  _T_3110_im = _RAND_5841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5842 = {1{`RANDOM}};
  _T_3111_re = _RAND_5842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5843 = {1{`RANDOM}};
  _T_3111_im = _RAND_5843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5844 = {1{`RANDOM}};
  _T_3112_re = _RAND_5844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5845 = {1{`RANDOM}};
  _T_3112_im = _RAND_5845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5846 = {1{`RANDOM}};
  _T_3113_re = _RAND_5846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5847 = {1{`RANDOM}};
  _T_3113_im = _RAND_5847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5848 = {1{`RANDOM}};
  _T_3114_re = _RAND_5848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5849 = {1{`RANDOM}};
  _T_3114_im = _RAND_5849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5850 = {1{`RANDOM}};
  _T_3115_re = _RAND_5850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5851 = {1{`RANDOM}};
  _T_3115_im = _RAND_5851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5852 = {1{`RANDOM}};
  _T_3116_re = _RAND_5852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5853 = {1{`RANDOM}};
  _T_3116_im = _RAND_5853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5854 = {1{`RANDOM}};
  _T_3117_re = _RAND_5854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5855 = {1{`RANDOM}};
  _T_3117_im = _RAND_5855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5856 = {1{`RANDOM}};
  _T_3118_re = _RAND_5856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5857 = {1{`RANDOM}};
  _T_3118_im = _RAND_5857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5858 = {1{`RANDOM}};
  _T_3119_re = _RAND_5858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5859 = {1{`RANDOM}};
  _T_3119_im = _RAND_5859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5860 = {1{`RANDOM}};
  _T_3120_re = _RAND_5860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5861 = {1{`RANDOM}};
  _T_3120_im = _RAND_5861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5862 = {1{`RANDOM}};
  _T_3121_re = _RAND_5862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5863 = {1{`RANDOM}};
  _T_3121_im = _RAND_5863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5864 = {1{`RANDOM}};
  _T_3122_re = _RAND_5864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5865 = {1{`RANDOM}};
  _T_3122_im = _RAND_5865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5866 = {1{`RANDOM}};
  _T_3123_re = _RAND_5866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5867 = {1{`RANDOM}};
  _T_3123_im = _RAND_5867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5868 = {1{`RANDOM}};
  _T_3124_re = _RAND_5868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5869 = {1{`RANDOM}};
  _T_3124_im = _RAND_5869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5870 = {1{`RANDOM}};
  _T_3125_re = _RAND_5870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5871 = {1{`RANDOM}};
  _T_3125_im = _RAND_5871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5872 = {1{`RANDOM}};
  _T_3126_re = _RAND_5872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5873 = {1{`RANDOM}};
  _T_3126_im = _RAND_5873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5874 = {1{`RANDOM}};
  _T_3127_re = _RAND_5874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5875 = {1{`RANDOM}};
  _T_3127_im = _RAND_5875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5876 = {1{`RANDOM}};
  _T_3128_re = _RAND_5876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5877 = {1{`RANDOM}};
  _T_3128_im = _RAND_5877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5878 = {1{`RANDOM}};
  _T_3129_re = _RAND_5878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5879 = {1{`RANDOM}};
  _T_3129_im = _RAND_5879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5880 = {1{`RANDOM}};
  _T_3130_re = _RAND_5880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5881 = {1{`RANDOM}};
  _T_3130_im = _RAND_5881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5882 = {1{`RANDOM}};
  _T_3131_re = _RAND_5882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5883 = {1{`RANDOM}};
  _T_3131_im = _RAND_5883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5884 = {1{`RANDOM}};
  _T_3132_re = _RAND_5884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5885 = {1{`RANDOM}};
  _T_3132_im = _RAND_5885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5886 = {1{`RANDOM}};
  _T_3133_re = _RAND_5886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5887 = {1{`RANDOM}};
  _T_3133_im = _RAND_5887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5888 = {1{`RANDOM}};
  _T_3134_re = _RAND_5888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5889 = {1{`RANDOM}};
  _T_3134_im = _RAND_5889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5890 = {1{`RANDOM}};
  _T_3135_re = _RAND_5890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5891 = {1{`RANDOM}};
  _T_3135_im = _RAND_5891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5892 = {1{`RANDOM}};
  _T_3136_re = _RAND_5892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5893 = {1{`RANDOM}};
  _T_3136_im = _RAND_5893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5894 = {1{`RANDOM}};
  _T_3137_re = _RAND_5894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5895 = {1{`RANDOM}};
  _T_3137_im = _RAND_5895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5896 = {1{`RANDOM}};
  _T_3138_re = _RAND_5896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5897 = {1{`RANDOM}};
  _T_3138_im = _RAND_5897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5898 = {1{`RANDOM}};
  _T_3139_re = _RAND_5898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5899 = {1{`RANDOM}};
  _T_3139_im = _RAND_5899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5900 = {1{`RANDOM}};
  _T_3140_re = _RAND_5900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5901 = {1{`RANDOM}};
  _T_3140_im = _RAND_5901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5902 = {1{`RANDOM}};
  _T_3141_re = _RAND_5902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5903 = {1{`RANDOM}};
  _T_3141_im = _RAND_5903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5904 = {1{`RANDOM}};
  _T_3142_re = _RAND_5904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5905 = {1{`RANDOM}};
  _T_3142_im = _RAND_5905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5906 = {1{`RANDOM}};
  _T_3143_re = _RAND_5906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5907 = {1{`RANDOM}};
  _T_3143_im = _RAND_5907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5908 = {1{`RANDOM}};
  _T_3144_re = _RAND_5908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5909 = {1{`RANDOM}};
  _T_3144_im = _RAND_5909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5910 = {1{`RANDOM}};
  _T_3145_re = _RAND_5910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5911 = {1{`RANDOM}};
  _T_3145_im = _RAND_5911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5912 = {1{`RANDOM}};
  _T_3146_re = _RAND_5912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5913 = {1{`RANDOM}};
  _T_3146_im = _RAND_5913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5914 = {1{`RANDOM}};
  _T_3147_re = _RAND_5914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5915 = {1{`RANDOM}};
  _T_3147_im = _RAND_5915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5916 = {1{`RANDOM}};
  _T_3148_re = _RAND_5916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5917 = {1{`RANDOM}};
  _T_3148_im = _RAND_5917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5918 = {1{`RANDOM}};
  _T_3149_re = _RAND_5918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5919 = {1{`RANDOM}};
  _T_3149_im = _RAND_5919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5920 = {1{`RANDOM}};
  _T_3150_re = _RAND_5920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5921 = {1{`RANDOM}};
  _T_3150_im = _RAND_5921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5922 = {1{`RANDOM}};
  _T_3151_re = _RAND_5922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5923 = {1{`RANDOM}};
  _T_3151_im = _RAND_5923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5924 = {1{`RANDOM}};
  _T_3152_re = _RAND_5924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5925 = {1{`RANDOM}};
  _T_3152_im = _RAND_5925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5926 = {1{`RANDOM}};
  _T_3153_re = _RAND_5926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5927 = {1{`RANDOM}};
  _T_3153_im = _RAND_5927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5928 = {1{`RANDOM}};
  _T_3154_re = _RAND_5928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5929 = {1{`RANDOM}};
  _T_3154_im = _RAND_5929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5930 = {1{`RANDOM}};
  _T_3155_re = _RAND_5930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5931 = {1{`RANDOM}};
  _T_3155_im = _RAND_5931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5932 = {1{`RANDOM}};
  _T_3156_re = _RAND_5932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5933 = {1{`RANDOM}};
  _T_3156_im = _RAND_5933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5934 = {1{`RANDOM}};
  _T_3157_re = _RAND_5934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5935 = {1{`RANDOM}};
  _T_3157_im = _RAND_5935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5936 = {1{`RANDOM}};
  _T_3158_re = _RAND_5936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5937 = {1{`RANDOM}};
  _T_3158_im = _RAND_5937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5938 = {1{`RANDOM}};
  _T_3159_re = _RAND_5938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5939 = {1{`RANDOM}};
  _T_3159_im = _RAND_5939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5940 = {1{`RANDOM}};
  _T_3160_re = _RAND_5940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5941 = {1{`RANDOM}};
  _T_3160_im = _RAND_5941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5942 = {1{`RANDOM}};
  _T_3161_re = _RAND_5942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5943 = {1{`RANDOM}};
  _T_3161_im = _RAND_5943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5944 = {1{`RANDOM}};
  _T_3162_re = _RAND_5944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5945 = {1{`RANDOM}};
  _T_3162_im = _RAND_5945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5946 = {1{`RANDOM}};
  _T_3163_re = _RAND_5946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5947 = {1{`RANDOM}};
  _T_3163_im = _RAND_5947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5948 = {1{`RANDOM}};
  _T_3164_re = _RAND_5948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5949 = {1{`RANDOM}};
  _T_3164_im = _RAND_5949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5950 = {1{`RANDOM}};
  _T_3165_re = _RAND_5950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5951 = {1{`RANDOM}};
  _T_3165_im = _RAND_5951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5952 = {1{`RANDOM}};
  _T_3166_re = _RAND_5952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5953 = {1{`RANDOM}};
  _T_3166_im = _RAND_5953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5954 = {1{`RANDOM}};
  _T_3167_re = _RAND_5954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5955 = {1{`RANDOM}};
  _T_3167_im = _RAND_5955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5956 = {1{`RANDOM}};
  _T_3168_re = _RAND_5956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5957 = {1{`RANDOM}};
  _T_3168_im = _RAND_5957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5958 = {1{`RANDOM}};
  _T_3169_re = _RAND_5958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5959 = {1{`RANDOM}};
  _T_3169_im = _RAND_5959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5960 = {1{`RANDOM}};
  _T_3170_re = _RAND_5960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5961 = {1{`RANDOM}};
  _T_3170_im = _RAND_5961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5962 = {1{`RANDOM}};
  _T_3171_re = _RAND_5962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5963 = {1{`RANDOM}};
  _T_3171_im = _RAND_5963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5964 = {1{`RANDOM}};
  _T_3172_re = _RAND_5964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5965 = {1{`RANDOM}};
  _T_3172_im = _RAND_5965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5966 = {1{`RANDOM}};
  _T_3173_re = _RAND_5966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5967 = {1{`RANDOM}};
  _T_3173_im = _RAND_5967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5968 = {1{`RANDOM}};
  _T_3174_re = _RAND_5968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5969 = {1{`RANDOM}};
  _T_3174_im = _RAND_5969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5970 = {1{`RANDOM}};
  _T_3175_re = _RAND_5970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5971 = {1{`RANDOM}};
  _T_3175_im = _RAND_5971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5972 = {1{`RANDOM}};
  _T_3176_re = _RAND_5972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5973 = {1{`RANDOM}};
  _T_3176_im = _RAND_5973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5974 = {1{`RANDOM}};
  _T_3177_re = _RAND_5974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5975 = {1{`RANDOM}};
  _T_3177_im = _RAND_5975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5976 = {1{`RANDOM}};
  _T_3178_re = _RAND_5976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5977 = {1{`RANDOM}};
  _T_3178_im = _RAND_5977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5978 = {1{`RANDOM}};
  _T_3179_re = _RAND_5978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5979 = {1{`RANDOM}};
  _T_3179_im = _RAND_5979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5980 = {1{`RANDOM}};
  _T_3180_re = _RAND_5980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5981 = {1{`RANDOM}};
  _T_3180_im = _RAND_5981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5982 = {1{`RANDOM}};
  _T_3181_re = _RAND_5982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5983 = {1{`RANDOM}};
  _T_3181_im = _RAND_5983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5984 = {1{`RANDOM}};
  _T_3182_re = _RAND_5984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5985 = {1{`RANDOM}};
  _T_3182_im = _RAND_5985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5986 = {1{`RANDOM}};
  _T_3183_re = _RAND_5986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5987 = {1{`RANDOM}};
  _T_3183_im = _RAND_5987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5988 = {1{`RANDOM}};
  _T_3184_re = _RAND_5988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5989 = {1{`RANDOM}};
  _T_3184_im = _RAND_5989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5990 = {1{`RANDOM}};
  _T_3185_re = _RAND_5990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5991 = {1{`RANDOM}};
  _T_3185_im = _RAND_5991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5992 = {1{`RANDOM}};
  _T_3186_re = _RAND_5992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5993 = {1{`RANDOM}};
  _T_3186_im = _RAND_5993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5994 = {1{`RANDOM}};
  _T_3187_re = _RAND_5994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5995 = {1{`RANDOM}};
  _T_3187_im = _RAND_5995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5996 = {1{`RANDOM}};
  _T_3188_re = _RAND_5996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5997 = {1{`RANDOM}};
  _T_3188_im = _RAND_5997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5998 = {1{`RANDOM}};
  _T_3189_re = _RAND_5998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5999 = {1{`RANDOM}};
  _T_3189_im = _RAND_5999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6000 = {1{`RANDOM}};
  _T_3190_re = _RAND_6000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6001 = {1{`RANDOM}};
  _T_3190_im = _RAND_6001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6002 = {1{`RANDOM}};
  _T_3191_re = _RAND_6002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6003 = {1{`RANDOM}};
  _T_3191_im = _RAND_6003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6004 = {1{`RANDOM}};
  _T_3192_re = _RAND_6004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6005 = {1{`RANDOM}};
  _T_3192_im = _RAND_6005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6006 = {1{`RANDOM}};
  _T_3193_re = _RAND_6006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6007 = {1{`RANDOM}};
  _T_3193_im = _RAND_6007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6008 = {1{`RANDOM}};
  _T_3194_re = _RAND_6008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6009 = {1{`RANDOM}};
  _T_3194_im = _RAND_6009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6010 = {1{`RANDOM}};
  _T_3195_re = _RAND_6010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6011 = {1{`RANDOM}};
  _T_3195_im = _RAND_6011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6012 = {1{`RANDOM}};
  _T_3196_re = _RAND_6012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6013 = {1{`RANDOM}};
  _T_3196_im = _RAND_6013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6014 = {1{`RANDOM}};
  _T_3197_re = _RAND_6014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6015 = {1{`RANDOM}};
  _T_3197_im = _RAND_6015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6016 = {1{`RANDOM}};
  _T_3198_re = _RAND_6016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6017 = {1{`RANDOM}};
  _T_3198_im = _RAND_6017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6018 = {1{`RANDOM}};
  _T_3199_re = _RAND_6018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6019 = {1{`RANDOM}};
  _T_3199_im = _RAND_6019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6020 = {1{`RANDOM}};
  _T_3200_re = _RAND_6020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6021 = {1{`RANDOM}};
  _T_3200_im = _RAND_6021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6022 = {1{`RANDOM}};
  _T_3201_re = _RAND_6022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6023 = {1{`RANDOM}};
  _T_3201_im = _RAND_6023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6024 = {1{`RANDOM}};
  _T_3202_re = _RAND_6024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6025 = {1{`RANDOM}};
  _T_3202_im = _RAND_6025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6026 = {1{`RANDOM}};
  _T_3203_re = _RAND_6026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6027 = {1{`RANDOM}};
  _T_3203_im = _RAND_6027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6028 = {1{`RANDOM}};
  _T_3204_re = _RAND_6028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6029 = {1{`RANDOM}};
  _T_3204_im = _RAND_6029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6030 = {1{`RANDOM}};
  _T_3205_re = _RAND_6030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6031 = {1{`RANDOM}};
  _T_3205_im = _RAND_6031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6032 = {1{`RANDOM}};
  _T_3206_re = _RAND_6032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6033 = {1{`RANDOM}};
  _T_3206_im = _RAND_6033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6034 = {1{`RANDOM}};
  _T_3207_re = _RAND_6034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6035 = {1{`RANDOM}};
  _T_3207_im = _RAND_6035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6036 = {1{`RANDOM}};
  _T_3208_re = _RAND_6036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6037 = {1{`RANDOM}};
  _T_3208_im = _RAND_6037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6038 = {1{`RANDOM}};
  _T_3209_re = _RAND_6038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6039 = {1{`RANDOM}};
  _T_3209_im = _RAND_6039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6040 = {1{`RANDOM}};
  _T_3210_re = _RAND_6040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6041 = {1{`RANDOM}};
  _T_3210_im = _RAND_6041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6042 = {1{`RANDOM}};
  _T_3211_re = _RAND_6042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6043 = {1{`RANDOM}};
  _T_3211_im = _RAND_6043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6044 = {1{`RANDOM}};
  _T_3212_re = _RAND_6044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6045 = {1{`RANDOM}};
  _T_3212_im = _RAND_6045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6046 = {1{`RANDOM}};
  _T_3213_re = _RAND_6046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6047 = {1{`RANDOM}};
  _T_3213_im = _RAND_6047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6048 = {1{`RANDOM}};
  _T_3214_re = _RAND_6048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6049 = {1{`RANDOM}};
  _T_3214_im = _RAND_6049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6050 = {1{`RANDOM}};
  _T_3215_re = _RAND_6050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6051 = {1{`RANDOM}};
  _T_3215_im = _RAND_6051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6052 = {1{`RANDOM}};
  _T_3216_re = _RAND_6052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6053 = {1{`RANDOM}};
  _T_3216_im = _RAND_6053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6054 = {1{`RANDOM}};
  _T_3217_re = _RAND_6054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6055 = {1{`RANDOM}};
  _T_3217_im = _RAND_6055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6056 = {1{`RANDOM}};
  _T_3218_re = _RAND_6056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6057 = {1{`RANDOM}};
  _T_3218_im = _RAND_6057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6058 = {1{`RANDOM}};
  _T_3219_re = _RAND_6058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6059 = {1{`RANDOM}};
  _T_3219_im = _RAND_6059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6060 = {1{`RANDOM}};
  _T_3220_re = _RAND_6060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6061 = {1{`RANDOM}};
  _T_3220_im = _RAND_6061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6062 = {1{`RANDOM}};
  _T_3221_re = _RAND_6062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6063 = {1{`RANDOM}};
  _T_3221_im = _RAND_6063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6064 = {1{`RANDOM}};
  _T_3222_re = _RAND_6064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6065 = {1{`RANDOM}};
  _T_3222_im = _RAND_6065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6066 = {1{`RANDOM}};
  _T_3223_re = _RAND_6066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6067 = {1{`RANDOM}};
  _T_3223_im = _RAND_6067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6068 = {1{`RANDOM}};
  _T_3224_re = _RAND_6068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6069 = {1{`RANDOM}};
  _T_3224_im = _RAND_6069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6070 = {1{`RANDOM}};
  _T_3225_re = _RAND_6070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6071 = {1{`RANDOM}};
  _T_3225_im = _RAND_6071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6072 = {1{`RANDOM}};
  _T_3226_re = _RAND_6072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6073 = {1{`RANDOM}};
  _T_3226_im = _RAND_6073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6074 = {1{`RANDOM}};
  _T_3227_re = _RAND_6074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6075 = {1{`RANDOM}};
  _T_3227_im = _RAND_6075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6076 = {1{`RANDOM}};
  _T_3228_re = _RAND_6076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6077 = {1{`RANDOM}};
  _T_3228_im = _RAND_6077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6078 = {1{`RANDOM}};
  _T_3229_re = _RAND_6078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6079 = {1{`RANDOM}};
  _T_3229_im = _RAND_6079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6080 = {1{`RANDOM}};
  _T_3230_re = _RAND_6080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6081 = {1{`RANDOM}};
  _T_3230_im = _RAND_6081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6082 = {1{`RANDOM}};
  _T_3231_re = _RAND_6082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6083 = {1{`RANDOM}};
  _T_3231_im = _RAND_6083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6084 = {1{`RANDOM}};
  _T_3232_re = _RAND_6084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6085 = {1{`RANDOM}};
  _T_3232_im = _RAND_6085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6086 = {1{`RANDOM}};
  _T_3233_re = _RAND_6086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6087 = {1{`RANDOM}};
  _T_3233_im = _RAND_6087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6088 = {1{`RANDOM}};
  _T_3234_re = _RAND_6088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6089 = {1{`RANDOM}};
  _T_3234_im = _RAND_6089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6090 = {1{`RANDOM}};
  _T_3235_re = _RAND_6090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6091 = {1{`RANDOM}};
  _T_3235_im = _RAND_6091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6092 = {1{`RANDOM}};
  _T_3236_re = _RAND_6092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6093 = {1{`RANDOM}};
  _T_3236_im = _RAND_6093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6094 = {1{`RANDOM}};
  _T_3237_re = _RAND_6094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6095 = {1{`RANDOM}};
  _T_3237_im = _RAND_6095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6096 = {1{`RANDOM}};
  _T_3238_re = _RAND_6096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6097 = {1{`RANDOM}};
  _T_3238_im = _RAND_6097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6098 = {1{`RANDOM}};
  _T_3239_re = _RAND_6098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6099 = {1{`RANDOM}};
  _T_3239_im = _RAND_6099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6100 = {1{`RANDOM}};
  _T_3240_re = _RAND_6100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6101 = {1{`RANDOM}};
  _T_3240_im = _RAND_6101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6102 = {1{`RANDOM}};
  _T_3241_re = _RAND_6102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6103 = {1{`RANDOM}};
  _T_3241_im = _RAND_6103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6104 = {1{`RANDOM}};
  _T_3242_re = _RAND_6104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6105 = {1{`RANDOM}};
  _T_3242_im = _RAND_6105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6106 = {1{`RANDOM}};
  _T_3243_re = _RAND_6106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6107 = {1{`RANDOM}};
  _T_3243_im = _RAND_6107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6108 = {1{`RANDOM}};
  _T_3244_re = _RAND_6108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6109 = {1{`RANDOM}};
  _T_3244_im = _RAND_6109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6110 = {1{`RANDOM}};
  _T_3245_re = _RAND_6110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6111 = {1{`RANDOM}};
  _T_3245_im = _RAND_6111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6112 = {1{`RANDOM}};
  _T_3246_re = _RAND_6112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6113 = {1{`RANDOM}};
  _T_3246_im = _RAND_6113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6114 = {1{`RANDOM}};
  _T_3247_re = _RAND_6114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6115 = {1{`RANDOM}};
  _T_3247_im = _RAND_6115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6116 = {1{`RANDOM}};
  _T_3248_re = _RAND_6116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6117 = {1{`RANDOM}};
  _T_3248_im = _RAND_6117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6118 = {1{`RANDOM}};
  _T_3249_re = _RAND_6118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6119 = {1{`RANDOM}};
  _T_3249_im = _RAND_6119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6120 = {1{`RANDOM}};
  _T_3250_re = _RAND_6120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6121 = {1{`RANDOM}};
  _T_3250_im = _RAND_6121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6122 = {1{`RANDOM}};
  _T_3251_re = _RAND_6122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6123 = {1{`RANDOM}};
  _T_3251_im = _RAND_6123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6124 = {1{`RANDOM}};
  _T_3252_re = _RAND_6124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6125 = {1{`RANDOM}};
  _T_3252_im = _RAND_6125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6126 = {1{`RANDOM}};
  _T_3253_re = _RAND_6126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6127 = {1{`RANDOM}};
  _T_3253_im = _RAND_6127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6128 = {1{`RANDOM}};
  _T_3254_re = _RAND_6128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6129 = {1{`RANDOM}};
  _T_3254_im = _RAND_6129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6130 = {1{`RANDOM}};
  _T_3255_re = _RAND_6130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6131 = {1{`RANDOM}};
  _T_3255_im = _RAND_6131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6132 = {1{`RANDOM}};
  _T_3256_re = _RAND_6132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6133 = {1{`RANDOM}};
  _T_3256_im = _RAND_6133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6134 = {1{`RANDOM}};
  _T_3257_re = _RAND_6134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6135 = {1{`RANDOM}};
  _T_3257_im = _RAND_6135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6136 = {1{`RANDOM}};
  _T_3258_re = _RAND_6136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6137 = {1{`RANDOM}};
  _T_3258_im = _RAND_6137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6138 = {1{`RANDOM}};
  _T_3259_re = _RAND_6138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6139 = {1{`RANDOM}};
  _T_3259_im = _RAND_6139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6140 = {1{`RANDOM}};
  _T_3260_re = _RAND_6140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6141 = {1{`RANDOM}};
  _T_3260_im = _RAND_6141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6142 = {1{`RANDOM}};
  _T_3261_re = _RAND_6142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6143 = {1{`RANDOM}};
  _T_3261_im = _RAND_6143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6144 = {1{`RANDOM}};
  _T_3262_re = _RAND_6144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6145 = {1{`RANDOM}};
  _T_3262_im = _RAND_6145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6146 = {1{`RANDOM}};
  _T_3268_re = _RAND_6146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6147 = {1{`RANDOM}};
  _T_3268_im = _RAND_6147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6148 = {1{`RANDOM}};
  _T_3269_re = _RAND_6148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6149 = {1{`RANDOM}};
  _T_3269_im = _RAND_6149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6150 = {1{`RANDOM}};
  _T_3270_re = _RAND_6150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6151 = {1{`RANDOM}};
  _T_3270_im = _RAND_6151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6152 = {1{`RANDOM}};
  _T_3271_re = _RAND_6152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6153 = {1{`RANDOM}};
  _T_3271_im = _RAND_6153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6154 = {1{`RANDOM}};
  _T_3272_re = _RAND_6154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6155 = {1{`RANDOM}};
  _T_3272_im = _RAND_6155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6156 = {1{`RANDOM}};
  _T_3273_re = _RAND_6156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6157 = {1{`RANDOM}};
  _T_3273_im = _RAND_6157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6158 = {1{`RANDOM}};
  _T_3274_re = _RAND_6158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6159 = {1{`RANDOM}};
  _T_3274_im = _RAND_6159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6160 = {1{`RANDOM}};
  _T_3275_re = _RAND_6160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6161 = {1{`RANDOM}};
  _T_3275_im = _RAND_6161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6162 = {1{`RANDOM}};
  _T_3276_re = _RAND_6162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6163 = {1{`RANDOM}};
  _T_3276_im = _RAND_6163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6164 = {1{`RANDOM}};
  _T_3277_re = _RAND_6164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6165 = {1{`RANDOM}};
  _T_3277_im = _RAND_6165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6166 = {1{`RANDOM}};
  _T_3278_re = _RAND_6166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6167 = {1{`RANDOM}};
  _T_3278_im = _RAND_6167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6168 = {1{`RANDOM}};
  _T_3279_re = _RAND_6168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6169 = {1{`RANDOM}};
  _T_3279_im = _RAND_6169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6170 = {1{`RANDOM}};
  _T_3280_re = _RAND_6170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6171 = {1{`RANDOM}};
  _T_3280_im = _RAND_6171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6172 = {1{`RANDOM}};
  _T_3281_re = _RAND_6172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6173 = {1{`RANDOM}};
  _T_3281_im = _RAND_6173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6174 = {1{`RANDOM}};
  _T_3282_re = _RAND_6174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6175 = {1{`RANDOM}};
  _T_3282_im = _RAND_6175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6176 = {1{`RANDOM}};
  _T_3283_re = _RAND_6176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6177 = {1{`RANDOM}};
  _T_3283_im = _RAND_6177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6178 = {1{`RANDOM}};
  _T_3284_re = _RAND_6178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6179 = {1{`RANDOM}};
  _T_3284_im = _RAND_6179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6180 = {1{`RANDOM}};
  _T_3285_re = _RAND_6180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6181 = {1{`RANDOM}};
  _T_3285_im = _RAND_6181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6182 = {1{`RANDOM}};
  _T_3286_re = _RAND_6182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6183 = {1{`RANDOM}};
  _T_3286_im = _RAND_6183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6184 = {1{`RANDOM}};
  _T_3287_re = _RAND_6184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6185 = {1{`RANDOM}};
  _T_3287_im = _RAND_6185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6186 = {1{`RANDOM}};
  _T_3288_re = _RAND_6186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6187 = {1{`RANDOM}};
  _T_3288_im = _RAND_6187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6188 = {1{`RANDOM}};
  _T_3289_re = _RAND_6188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6189 = {1{`RANDOM}};
  _T_3289_im = _RAND_6189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6190 = {1{`RANDOM}};
  _T_3290_re = _RAND_6190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6191 = {1{`RANDOM}};
  _T_3290_im = _RAND_6191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6192 = {1{`RANDOM}};
  _T_3291_re = _RAND_6192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6193 = {1{`RANDOM}};
  _T_3291_im = _RAND_6193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6194 = {1{`RANDOM}};
  _T_3292_re = _RAND_6194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6195 = {1{`RANDOM}};
  _T_3292_im = _RAND_6195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6196 = {1{`RANDOM}};
  _T_3293_re = _RAND_6196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6197 = {1{`RANDOM}};
  _T_3293_im = _RAND_6197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6198 = {1{`RANDOM}};
  _T_3294_re = _RAND_6198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6199 = {1{`RANDOM}};
  _T_3294_im = _RAND_6199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6200 = {1{`RANDOM}};
  _T_3295_re = _RAND_6200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6201 = {1{`RANDOM}};
  _T_3295_im = _RAND_6201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6202 = {1{`RANDOM}};
  _T_3296_re = _RAND_6202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6203 = {1{`RANDOM}};
  _T_3296_im = _RAND_6203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6204 = {1{`RANDOM}};
  _T_3297_re = _RAND_6204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6205 = {1{`RANDOM}};
  _T_3297_im = _RAND_6205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6206 = {1{`RANDOM}};
  _T_3298_re = _RAND_6206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6207 = {1{`RANDOM}};
  _T_3298_im = _RAND_6207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6208 = {1{`RANDOM}};
  _T_3299_re = _RAND_6208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6209 = {1{`RANDOM}};
  _T_3299_im = _RAND_6209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6210 = {1{`RANDOM}};
  _T_3300_re = _RAND_6210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6211 = {1{`RANDOM}};
  _T_3300_im = _RAND_6211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6212 = {1{`RANDOM}};
  _T_3301_re = _RAND_6212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6213 = {1{`RANDOM}};
  _T_3301_im = _RAND_6213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6214 = {1{`RANDOM}};
  _T_3302_re = _RAND_6214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6215 = {1{`RANDOM}};
  _T_3302_im = _RAND_6215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6216 = {1{`RANDOM}};
  _T_3303_re = _RAND_6216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6217 = {1{`RANDOM}};
  _T_3303_im = _RAND_6217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6218 = {1{`RANDOM}};
  _T_3304_re = _RAND_6218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6219 = {1{`RANDOM}};
  _T_3304_im = _RAND_6219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6220 = {1{`RANDOM}};
  _T_3305_re = _RAND_6220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6221 = {1{`RANDOM}};
  _T_3305_im = _RAND_6221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6222 = {1{`RANDOM}};
  _T_3306_re = _RAND_6222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6223 = {1{`RANDOM}};
  _T_3306_im = _RAND_6223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6224 = {1{`RANDOM}};
  _T_3307_re = _RAND_6224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6225 = {1{`RANDOM}};
  _T_3307_im = _RAND_6225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6226 = {1{`RANDOM}};
  _T_3308_re = _RAND_6226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6227 = {1{`RANDOM}};
  _T_3308_im = _RAND_6227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6228 = {1{`RANDOM}};
  _T_3309_re = _RAND_6228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6229 = {1{`RANDOM}};
  _T_3309_im = _RAND_6229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6230 = {1{`RANDOM}};
  _T_3310_re = _RAND_6230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6231 = {1{`RANDOM}};
  _T_3310_im = _RAND_6231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6232 = {1{`RANDOM}};
  _T_3311_re = _RAND_6232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6233 = {1{`RANDOM}};
  _T_3311_im = _RAND_6233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6234 = {1{`RANDOM}};
  _T_3312_re = _RAND_6234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6235 = {1{`RANDOM}};
  _T_3312_im = _RAND_6235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6236 = {1{`RANDOM}};
  _T_3313_re = _RAND_6236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6237 = {1{`RANDOM}};
  _T_3313_im = _RAND_6237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6238 = {1{`RANDOM}};
  _T_3314_re = _RAND_6238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6239 = {1{`RANDOM}};
  _T_3314_im = _RAND_6239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6240 = {1{`RANDOM}};
  _T_3315_re = _RAND_6240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6241 = {1{`RANDOM}};
  _T_3315_im = _RAND_6241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6242 = {1{`RANDOM}};
  _T_3316_re = _RAND_6242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6243 = {1{`RANDOM}};
  _T_3316_im = _RAND_6243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6244 = {1{`RANDOM}};
  _T_3317_re = _RAND_6244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6245 = {1{`RANDOM}};
  _T_3317_im = _RAND_6245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6246 = {1{`RANDOM}};
  _T_3318_re = _RAND_6246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6247 = {1{`RANDOM}};
  _T_3318_im = _RAND_6247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6248 = {1{`RANDOM}};
  _T_3319_re = _RAND_6248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6249 = {1{`RANDOM}};
  _T_3319_im = _RAND_6249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6250 = {1{`RANDOM}};
  _T_3320_re = _RAND_6250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6251 = {1{`RANDOM}};
  _T_3320_im = _RAND_6251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6252 = {1{`RANDOM}};
  _T_3321_re = _RAND_6252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6253 = {1{`RANDOM}};
  _T_3321_im = _RAND_6253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6254 = {1{`RANDOM}};
  _T_3322_re = _RAND_6254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6255 = {1{`RANDOM}};
  _T_3322_im = _RAND_6255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6256 = {1{`RANDOM}};
  _T_3323_re = _RAND_6256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6257 = {1{`RANDOM}};
  _T_3323_im = _RAND_6257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6258 = {1{`RANDOM}};
  _T_3324_re = _RAND_6258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6259 = {1{`RANDOM}};
  _T_3324_im = _RAND_6259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6260 = {1{`RANDOM}};
  _T_3325_re = _RAND_6260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6261 = {1{`RANDOM}};
  _T_3325_im = _RAND_6261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6262 = {1{`RANDOM}};
  _T_3326_re = _RAND_6262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6263 = {1{`RANDOM}};
  _T_3326_im = _RAND_6263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6264 = {1{`RANDOM}};
  _T_3327_re = _RAND_6264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6265 = {1{`RANDOM}};
  _T_3327_im = _RAND_6265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6266 = {1{`RANDOM}};
  _T_3328_re = _RAND_6266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6267 = {1{`RANDOM}};
  _T_3328_im = _RAND_6267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6268 = {1{`RANDOM}};
  _T_3329_re = _RAND_6268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6269 = {1{`RANDOM}};
  _T_3329_im = _RAND_6269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6270 = {1{`RANDOM}};
  _T_3330_re = _RAND_6270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6271 = {1{`RANDOM}};
  _T_3330_im = _RAND_6271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6272 = {1{`RANDOM}};
  _T_3331_re = _RAND_6272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6273 = {1{`RANDOM}};
  _T_3331_im = _RAND_6273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6274 = {1{`RANDOM}};
  _T_3332_re = _RAND_6274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6275 = {1{`RANDOM}};
  _T_3332_im = _RAND_6275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6276 = {1{`RANDOM}};
  _T_3333_re = _RAND_6276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6277 = {1{`RANDOM}};
  _T_3333_im = _RAND_6277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6278 = {1{`RANDOM}};
  _T_3334_re = _RAND_6278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6279 = {1{`RANDOM}};
  _T_3334_im = _RAND_6279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6280 = {1{`RANDOM}};
  _T_3335_re = _RAND_6280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6281 = {1{`RANDOM}};
  _T_3335_im = _RAND_6281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6282 = {1{`RANDOM}};
  _T_3336_re = _RAND_6282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6283 = {1{`RANDOM}};
  _T_3336_im = _RAND_6283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6284 = {1{`RANDOM}};
  _T_3337_re = _RAND_6284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6285 = {1{`RANDOM}};
  _T_3337_im = _RAND_6285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6286 = {1{`RANDOM}};
  _T_3338_re = _RAND_6286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6287 = {1{`RANDOM}};
  _T_3338_im = _RAND_6287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6288 = {1{`RANDOM}};
  _T_3339_re = _RAND_6288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6289 = {1{`RANDOM}};
  _T_3339_im = _RAND_6289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6290 = {1{`RANDOM}};
  _T_3340_re = _RAND_6290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6291 = {1{`RANDOM}};
  _T_3340_im = _RAND_6291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6292 = {1{`RANDOM}};
  _T_3341_re = _RAND_6292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6293 = {1{`RANDOM}};
  _T_3341_im = _RAND_6293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6294 = {1{`RANDOM}};
  _T_3342_re = _RAND_6294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6295 = {1{`RANDOM}};
  _T_3342_im = _RAND_6295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6296 = {1{`RANDOM}};
  _T_3343_re = _RAND_6296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6297 = {1{`RANDOM}};
  _T_3343_im = _RAND_6297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6298 = {1{`RANDOM}};
  _T_3344_re = _RAND_6298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6299 = {1{`RANDOM}};
  _T_3344_im = _RAND_6299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6300 = {1{`RANDOM}};
  _T_3345_re = _RAND_6300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6301 = {1{`RANDOM}};
  _T_3345_im = _RAND_6301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6302 = {1{`RANDOM}};
  _T_3346_re = _RAND_6302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6303 = {1{`RANDOM}};
  _T_3346_im = _RAND_6303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6304 = {1{`RANDOM}};
  _T_3347_re = _RAND_6304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6305 = {1{`RANDOM}};
  _T_3347_im = _RAND_6305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6306 = {1{`RANDOM}};
  _T_3348_re = _RAND_6306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6307 = {1{`RANDOM}};
  _T_3348_im = _RAND_6307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6308 = {1{`RANDOM}};
  _T_3349_re = _RAND_6308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6309 = {1{`RANDOM}};
  _T_3349_im = _RAND_6309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6310 = {1{`RANDOM}};
  _T_3350_re = _RAND_6310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6311 = {1{`RANDOM}};
  _T_3350_im = _RAND_6311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6312 = {1{`RANDOM}};
  _T_3351_re = _RAND_6312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6313 = {1{`RANDOM}};
  _T_3351_im = _RAND_6313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6314 = {1{`RANDOM}};
  _T_3352_re = _RAND_6314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6315 = {1{`RANDOM}};
  _T_3352_im = _RAND_6315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6316 = {1{`RANDOM}};
  _T_3353_re = _RAND_6316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6317 = {1{`RANDOM}};
  _T_3353_im = _RAND_6317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6318 = {1{`RANDOM}};
  _T_3354_re = _RAND_6318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6319 = {1{`RANDOM}};
  _T_3354_im = _RAND_6319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6320 = {1{`RANDOM}};
  _T_3355_re = _RAND_6320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6321 = {1{`RANDOM}};
  _T_3355_im = _RAND_6321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6322 = {1{`RANDOM}};
  _T_3356_re = _RAND_6322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6323 = {1{`RANDOM}};
  _T_3356_im = _RAND_6323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6324 = {1{`RANDOM}};
  _T_3357_re = _RAND_6324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6325 = {1{`RANDOM}};
  _T_3357_im = _RAND_6325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6326 = {1{`RANDOM}};
  _T_3358_re = _RAND_6326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6327 = {1{`RANDOM}};
  _T_3358_im = _RAND_6327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6328 = {1{`RANDOM}};
  _T_3359_re = _RAND_6328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6329 = {1{`RANDOM}};
  _T_3359_im = _RAND_6329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6330 = {1{`RANDOM}};
  _T_3360_re = _RAND_6330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6331 = {1{`RANDOM}};
  _T_3360_im = _RAND_6331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6332 = {1{`RANDOM}};
  _T_3361_re = _RAND_6332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6333 = {1{`RANDOM}};
  _T_3361_im = _RAND_6333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6334 = {1{`RANDOM}};
  _T_3362_re = _RAND_6334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6335 = {1{`RANDOM}};
  _T_3362_im = _RAND_6335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6336 = {1{`RANDOM}};
  _T_3363_re = _RAND_6336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6337 = {1{`RANDOM}};
  _T_3363_im = _RAND_6337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6338 = {1{`RANDOM}};
  _T_3364_re = _RAND_6338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6339 = {1{`RANDOM}};
  _T_3364_im = _RAND_6339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6340 = {1{`RANDOM}};
  _T_3365_re = _RAND_6340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6341 = {1{`RANDOM}};
  _T_3365_im = _RAND_6341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6342 = {1{`RANDOM}};
  _T_3366_re = _RAND_6342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6343 = {1{`RANDOM}};
  _T_3366_im = _RAND_6343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6344 = {1{`RANDOM}};
  _T_3367_re = _RAND_6344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6345 = {1{`RANDOM}};
  _T_3367_im = _RAND_6345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6346 = {1{`RANDOM}};
  _T_3368_re = _RAND_6346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6347 = {1{`RANDOM}};
  _T_3368_im = _RAND_6347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6348 = {1{`RANDOM}};
  _T_3369_re = _RAND_6348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6349 = {1{`RANDOM}};
  _T_3369_im = _RAND_6349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6350 = {1{`RANDOM}};
  _T_3370_re = _RAND_6350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6351 = {1{`RANDOM}};
  _T_3370_im = _RAND_6351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6352 = {1{`RANDOM}};
  _T_3371_re = _RAND_6352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6353 = {1{`RANDOM}};
  _T_3371_im = _RAND_6353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6354 = {1{`RANDOM}};
  _T_3372_re = _RAND_6354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6355 = {1{`RANDOM}};
  _T_3372_im = _RAND_6355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6356 = {1{`RANDOM}};
  _T_3373_re = _RAND_6356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6357 = {1{`RANDOM}};
  _T_3373_im = _RAND_6357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6358 = {1{`RANDOM}};
  _T_3374_re = _RAND_6358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6359 = {1{`RANDOM}};
  _T_3374_im = _RAND_6359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6360 = {1{`RANDOM}};
  _T_3375_re = _RAND_6360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6361 = {1{`RANDOM}};
  _T_3375_im = _RAND_6361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6362 = {1{`RANDOM}};
  _T_3376_re = _RAND_6362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6363 = {1{`RANDOM}};
  _T_3376_im = _RAND_6363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6364 = {1{`RANDOM}};
  _T_3377_re = _RAND_6364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6365 = {1{`RANDOM}};
  _T_3377_im = _RAND_6365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6366 = {1{`RANDOM}};
  _T_3378_re = _RAND_6366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6367 = {1{`RANDOM}};
  _T_3378_im = _RAND_6367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6368 = {1{`RANDOM}};
  _T_3379_re = _RAND_6368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6369 = {1{`RANDOM}};
  _T_3379_im = _RAND_6369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6370 = {1{`RANDOM}};
  _T_3380_re = _RAND_6370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6371 = {1{`RANDOM}};
  _T_3380_im = _RAND_6371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6372 = {1{`RANDOM}};
  _T_3381_re = _RAND_6372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6373 = {1{`RANDOM}};
  _T_3381_im = _RAND_6373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6374 = {1{`RANDOM}};
  _T_3382_re = _RAND_6374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6375 = {1{`RANDOM}};
  _T_3382_im = _RAND_6375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6376 = {1{`RANDOM}};
  _T_3383_re = _RAND_6376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6377 = {1{`RANDOM}};
  _T_3383_im = _RAND_6377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6378 = {1{`RANDOM}};
  _T_3384_re = _RAND_6378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6379 = {1{`RANDOM}};
  _T_3384_im = _RAND_6379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6380 = {1{`RANDOM}};
  _T_3385_re = _RAND_6380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6381 = {1{`RANDOM}};
  _T_3385_im = _RAND_6381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6382 = {1{`RANDOM}};
  _T_3386_re = _RAND_6382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6383 = {1{`RANDOM}};
  _T_3386_im = _RAND_6383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6384 = {1{`RANDOM}};
  _T_3387_re = _RAND_6384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6385 = {1{`RANDOM}};
  _T_3387_im = _RAND_6385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6386 = {1{`RANDOM}};
  _T_3388_re = _RAND_6386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6387 = {1{`RANDOM}};
  _T_3388_im = _RAND_6387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6388 = {1{`RANDOM}};
  _T_3389_re = _RAND_6388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6389 = {1{`RANDOM}};
  _T_3389_im = _RAND_6389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6390 = {1{`RANDOM}};
  _T_3390_re = _RAND_6390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6391 = {1{`RANDOM}};
  _T_3390_im = _RAND_6391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6392 = {1{`RANDOM}};
  _T_3391_re = _RAND_6392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6393 = {1{`RANDOM}};
  _T_3391_im = _RAND_6393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6394 = {1{`RANDOM}};
  _T_3392_re = _RAND_6394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6395 = {1{`RANDOM}};
  _T_3392_im = _RAND_6395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6396 = {1{`RANDOM}};
  _T_3393_re = _RAND_6396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6397 = {1{`RANDOM}};
  _T_3393_im = _RAND_6397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6398 = {1{`RANDOM}};
  _T_3394_re = _RAND_6398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6399 = {1{`RANDOM}};
  _T_3394_im = _RAND_6399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6400 = {1{`RANDOM}};
  _T_3395_re = _RAND_6400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6401 = {1{`RANDOM}};
  _T_3395_im = _RAND_6401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6402 = {1{`RANDOM}};
  _T_3396_re = _RAND_6402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6403 = {1{`RANDOM}};
  _T_3396_im = _RAND_6403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6404 = {1{`RANDOM}};
  _T_3397_re = _RAND_6404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6405 = {1{`RANDOM}};
  _T_3397_im = _RAND_6405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6406 = {1{`RANDOM}};
  _T_3398_re = _RAND_6406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6407 = {1{`RANDOM}};
  _T_3398_im = _RAND_6407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6408 = {1{`RANDOM}};
  _T_3399_re = _RAND_6408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6409 = {1{`RANDOM}};
  _T_3399_im = _RAND_6409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6410 = {1{`RANDOM}};
  _T_3400_re = _RAND_6410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6411 = {1{`RANDOM}};
  _T_3400_im = _RAND_6411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6412 = {1{`RANDOM}};
  _T_3401_re = _RAND_6412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6413 = {1{`RANDOM}};
  _T_3401_im = _RAND_6413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6414 = {1{`RANDOM}};
  _T_3402_re = _RAND_6414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6415 = {1{`RANDOM}};
  _T_3402_im = _RAND_6415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6416 = {1{`RANDOM}};
  _T_3403_re = _RAND_6416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6417 = {1{`RANDOM}};
  _T_3403_im = _RAND_6417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6418 = {1{`RANDOM}};
  _T_3404_re = _RAND_6418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6419 = {1{`RANDOM}};
  _T_3404_im = _RAND_6419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6420 = {1{`RANDOM}};
  _T_3405_re = _RAND_6420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6421 = {1{`RANDOM}};
  _T_3405_im = _RAND_6421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6422 = {1{`RANDOM}};
  _T_3406_re = _RAND_6422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6423 = {1{`RANDOM}};
  _T_3406_im = _RAND_6423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6424 = {1{`RANDOM}};
  _T_3407_re = _RAND_6424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6425 = {1{`RANDOM}};
  _T_3407_im = _RAND_6425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6426 = {1{`RANDOM}};
  _T_3408_re = _RAND_6426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6427 = {1{`RANDOM}};
  _T_3408_im = _RAND_6427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6428 = {1{`RANDOM}};
  _T_3409_re = _RAND_6428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6429 = {1{`RANDOM}};
  _T_3409_im = _RAND_6429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6430 = {1{`RANDOM}};
  _T_3410_re = _RAND_6430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6431 = {1{`RANDOM}};
  _T_3410_im = _RAND_6431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6432 = {1{`RANDOM}};
  _T_3411_re = _RAND_6432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6433 = {1{`RANDOM}};
  _T_3411_im = _RAND_6433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6434 = {1{`RANDOM}};
  _T_3412_re = _RAND_6434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6435 = {1{`RANDOM}};
  _T_3412_im = _RAND_6435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6436 = {1{`RANDOM}};
  _T_3413_re = _RAND_6436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6437 = {1{`RANDOM}};
  _T_3413_im = _RAND_6437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6438 = {1{`RANDOM}};
  _T_3414_re = _RAND_6438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6439 = {1{`RANDOM}};
  _T_3414_im = _RAND_6439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6440 = {1{`RANDOM}};
  _T_3415_re = _RAND_6440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6441 = {1{`RANDOM}};
  _T_3415_im = _RAND_6441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6442 = {1{`RANDOM}};
  _T_3416_re = _RAND_6442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6443 = {1{`RANDOM}};
  _T_3416_im = _RAND_6443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6444 = {1{`RANDOM}};
  _T_3417_re = _RAND_6444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6445 = {1{`RANDOM}};
  _T_3417_im = _RAND_6445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6446 = {1{`RANDOM}};
  _T_3418_re = _RAND_6446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6447 = {1{`RANDOM}};
  _T_3418_im = _RAND_6447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6448 = {1{`RANDOM}};
  _T_3419_re = _RAND_6448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6449 = {1{`RANDOM}};
  _T_3419_im = _RAND_6449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6450 = {1{`RANDOM}};
  _T_3420_re = _RAND_6450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6451 = {1{`RANDOM}};
  _T_3420_im = _RAND_6451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6452 = {1{`RANDOM}};
  _T_3421_re = _RAND_6452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6453 = {1{`RANDOM}};
  _T_3421_im = _RAND_6453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6454 = {1{`RANDOM}};
  _T_3422_re = _RAND_6454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6455 = {1{`RANDOM}};
  _T_3422_im = _RAND_6455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6456 = {1{`RANDOM}};
  _T_3423_re = _RAND_6456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6457 = {1{`RANDOM}};
  _T_3423_im = _RAND_6457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6458 = {1{`RANDOM}};
  _T_3424_re = _RAND_6458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6459 = {1{`RANDOM}};
  _T_3424_im = _RAND_6459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6460 = {1{`RANDOM}};
  _T_3425_re = _RAND_6460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6461 = {1{`RANDOM}};
  _T_3425_im = _RAND_6461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6462 = {1{`RANDOM}};
  _T_3426_re = _RAND_6462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6463 = {1{`RANDOM}};
  _T_3426_im = _RAND_6463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6464 = {1{`RANDOM}};
  _T_3427_re = _RAND_6464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6465 = {1{`RANDOM}};
  _T_3427_im = _RAND_6465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6466 = {1{`RANDOM}};
  _T_3428_re = _RAND_6466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6467 = {1{`RANDOM}};
  _T_3428_im = _RAND_6467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6468 = {1{`RANDOM}};
  _T_3429_re = _RAND_6468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6469 = {1{`RANDOM}};
  _T_3429_im = _RAND_6469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6470 = {1{`RANDOM}};
  _T_3430_re = _RAND_6470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6471 = {1{`RANDOM}};
  _T_3430_im = _RAND_6471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6472 = {1{`RANDOM}};
  _T_3431_re = _RAND_6472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6473 = {1{`RANDOM}};
  _T_3431_im = _RAND_6473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6474 = {1{`RANDOM}};
  _T_3432_re = _RAND_6474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6475 = {1{`RANDOM}};
  _T_3432_im = _RAND_6475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6476 = {1{`RANDOM}};
  _T_3433_re = _RAND_6476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6477 = {1{`RANDOM}};
  _T_3433_im = _RAND_6477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6478 = {1{`RANDOM}};
  _T_3434_re = _RAND_6478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6479 = {1{`RANDOM}};
  _T_3434_im = _RAND_6479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6480 = {1{`RANDOM}};
  _T_3435_re = _RAND_6480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6481 = {1{`RANDOM}};
  _T_3435_im = _RAND_6481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6482 = {1{`RANDOM}};
  _T_3436_re = _RAND_6482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6483 = {1{`RANDOM}};
  _T_3436_im = _RAND_6483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6484 = {1{`RANDOM}};
  _T_3437_re = _RAND_6484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6485 = {1{`RANDOM}};
  _T_3437_im = _RAND_6485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6486 = {1{`RANDOM}};
  _T_3438_re = _RAND_6486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6487 = {1{`RANDOM}};
  _T_3438_im = _RAND_6487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6488 = {1{`RANDOM}};
  _T_3439_re = _RAND_6488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6489 = {1{`RANDOM}};
  _T_3439_im = _RAND_6489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6490 = {1{`RANDOM}};
  _T_3440_re = _RAND_6490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6491 = {1{`RANDOM}};
  _T_3440_im = _RAND_6491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6492 = {1{`RANDOM}};
  _T_3441_re = _RAND_6492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6493 = {1{`RANDOM}};
  _T_3441_im = _RAND_6493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6494 = {1{`RANDOM}};
  _T_3442_re = _RAND_6494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6495 = {1{`RANDOM}};
  _T_3442_im = _RAND_6495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6496 = {1{`RANDOM}};
  _T_3443_re = _RAND_6496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6497 = {1{`RANDOM}};
  _T_3443_im = _RAND_6497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6498 = {1{`RANDOM}};
  _T_3444_re = _RAND_6498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6499 = {1{`RANDOM}};
  _T_3444_im = _RAND_6499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6500 = {1{`RANDOM}};
  _T_3445_re = _RAND_6500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6501 = {1{`RANDOM}};
  _T_3445_im = _RAND_6501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6502 = {1{`RANDOM}};
  _T_3446_re = _RAND_6502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6503 = {1{`RANDOM}};
  _T_3446_im = _RAND_6503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6504 = {1{`RANDOM}};
  _T_3447_re = _RAND_6504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6505 = {1{`RANDOM}};
  _T_3447_im = _RAND_6505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6506 = {1{`RANDOM}};
  _T_3448_re = _RAND_6506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6507 = {1{`RANDOM}};
  _T_3448_im = _RAND_6507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6508 = {1{`RANDOM}};
  _T_3449_re = _RAND_6508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6509 = {1{`RANDOM}};
  _T_3449_im = _RAND_6509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6510 = {1{`RANDOM}};
  _T_3450_re = _RAND_6510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6511 = {1{`RANDOM}};
  _T_3450_im = _RAND_6511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6512 = {1{`RANDOM}};
  _T_3451_re = _RAND_6512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6513 = {1{`RANDOM}};
  _T_3451_im = _RAND_6513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6514 = {1{`RANDOM}};
  _T_3452_re = _RAND_6514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6515 = {1{`RANDOM}};
  _T_3452_im = _RAND_6515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6516 = {1{`RANDOM}};
  _T_3453_re = _RAND_6516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6517 = {1{`RANDOM}};
  _T_3453_im = _RAND_6517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6518 = {1{`RANDOM}};
  _T_3454_re = _RAND_6518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6519 = {1{`RANDOM}};
  _T_3454_im = _RAND_6519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6520 = {1{`RANDOM}};
  _T_3455_re = _RAND_6520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6521 = {1{`RANDOM}};
  _T_3455_im = _RAND_6521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6522 = {1{`RANDOM}};
  _T_3456_re = _RAND_6522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6523 = {1{`RANDOM}};
  _T_3456_im = _RAND_6523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6524 = {1{`RANDOM}};
  _T_3457_re = _RAND_6524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6525 = {1{`RANDOM}};
  _T_3457_im = _RAND_6525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6526 = {1{`RANDOM}};
  _T_3458_re = _RAND_6526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6527 = {1{`RANDOM}};
  _T_3458_im = _RAND_6527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6528 = {1{`RANDOM}};
  _T_3459_re = _RAND_6528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6529 = {1{`RANDOM}};
  _T_3459_im = _RAND_6529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6530 = {1{`RANDOM}};
  _T_3460_re = _RAND_6530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6531 = {1{`RANDOM}};
  _T_3460_im = _RAND_6531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6532 = {1{`RANDOM}};
  _T_3461_re = _RAND_6532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6533 = {1{`RANDOM}};
  _T_3461_im = _RAND_6533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6534 = {1{`RANDOM}};
  _T_3462_re = _RAND_6534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6535 = {1{`RANDOM}};
  _T_3462_im = _RAND_6535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6536 = {1{`RANDOM}};
  _T_3463_re = _RAND_6536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6537 = {1{`RANDOM}};
  _T_3463_im = _RAND_6537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6538 = {1{`RANDOM}};
  _T_3464_re = _RAND_6538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6539 = {1{`RANDOM}};
  _T_3464_im = _RAND_6539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6540 = {1{`RANDOM}};
  _T_3465_re = _RAND_6540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6541 = {1{`RANDOM}};
  _T_3465_im = _RAND_6541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6542 = {1{`RANDOM}};
  _T_3466_re = _RAND_6542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6543 = {1{`RANDOM}};
  _T_3466_im = _RAND_6543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6544 = {1{`RANDOM}};
  _T_3467_re = _RAND_6544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6545 = {1{`RANDOM}};
  _T_3467_im = _RAND_6545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6546 = {1{`RANDOM}};
  _T_3468_re = _RAND_6546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6547 = {1{`RANDOM}};
  _T_3468_im = _RAND_6547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6548 = {1{`RANDOM}};
  _T_3469_re = _RAND_6548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6549 = {1{`RANDOM}};
  _T_3469_im = _RAND_6549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6550 = {1{`RANDOM}};
  _T_3470_re = _RAND_6550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6551 = {1{`RANDOM}};
  _T_3470_im = _RAND_6551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6552 = {1{`RANDOM}};
  _T_3471_re = _RAND_6552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6553 = {1{`RANDOM}};
  _T_3471_im = _RAND_6553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6554 = {1{`RANDOM}};
  _T_3472_re = _RAND_6554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6555 = {1{`RANDOM}};
  _T_3472_im = _RAND_6555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6556 = {1{`RANDOM}};
  _T_3473_re = _RAND_6556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6557 = {1{`RANDOM}};
  _T_3473_im = _RAND_6557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6558 = {1{`RANDOM}};
  _T_3474_re = _RAND_6558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6559 = {1{`RANDOM}};
  _T_3474_im = _RAND_6559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6560 = {1{`RANDOM}};
  _T_3475_re = _RAND_6560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6561 = {1{`RANDOM}};
  _T_3475_im = _RAND_6561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6562 = {1{`RANDOM}};
  _T_3476_re = _RAND_6562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6563 = {1{`RANDOM}};
  _T_3476_im = _RAND_6563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6564 = {1{`RANDOM}};
  _T_3477_re = _RAND_6564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6565 = {1{`RANDOM}};
  _T_3477_im = _RAND_6565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6566 = {1{`RANDOM}};
  _T_3478_re = _RAND_6566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6567 = {1{`RANDOM}};
  _T_3478_im = _RAND_6567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6568 = {1{`RANDOM}};
  _T_3479_re = _RAND_6568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6569 = {1{`RANDOM}};
  _T_3479_im = _RAND_6569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6570 = {1{`RANDOM}};
  _T_3480_re = _RAND_6570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6571 = {1{`RANDOM}};
  _T_3480_im = _RAND_6571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6572 = {1{`RANDOM}};
  _T_3481_re = _RAND_6572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6573 = {1{`RANDOM}};
  _T_3481_im = _RAND_6573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6574 = {1{`RANDOM}};
  _T_3482_re = _RAND_6574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6575 = {1{`RANDOM}};
  _T_3482_im = _RAND_6575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6576 = {1{`RANDOM}};
  _T_3483_re = _RAND_6576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6577 = {1{`RANDOM}};
  _T_3483_im = _RAND_6577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6578 = {1{`RANDOM}};
  _T_3484_re = _RAND_6578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6579 = {1{`RANDOM}};
  _T_3484_im = _RAND_6579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6580 = {1{`RANDOM}};
  _T_3485_re = _RAND_6580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6581 = {1{`RANDOM}};
  _T_3485_im = _RAND_6581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6582 = {1{`RANDOM}};
  _T_3486_re = _RAND_6582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6583 = {1{`RANDOM}};
  _T_3486_im = _RAND_6583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6584 = {1{`RANDOM}};
  _T_3487_re = _RAND_6584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6585 = {1{`RANDOM}};
  _T_3487_im = _RAND_6585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6586 = {1{`RANDOM}};
  _T_3488_re = _RAND_6586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6587 = {1{`RANDOM}};
  _T_3488_im = _RAND_6587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6588 = {1{`RANDOM}};
  _T_3489_re = _RAND_6588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6589 = {1{`RANDOM}};
  _T_3489_im = _RAND_6589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6590 = {1{`RANDOM}};
  _T_3490_re = _RAND_6590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6591 = {1{`RANDOM}};
  _T_3490_im = _RAND_6591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6592 = {1{`RANDOM}};
  _T_3491_re = _RAND_6592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6593 = {1{`RANDOM}};
  _T_3491_im = _RAND_6593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6594 = {1{`RANDOM}};
  _T_3492_re = _RAND_6594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6595 = {1{`RANDOM}};
  _T_3492_im = _RAND_6595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6596 = {1{`RANDOM}};
  _T_3493_re = _RAND_6596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6597 = {1{`RANDOM}};
  _T_3493_im = _RAND_6597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6598 = {1{`RANDOM}};
  _T_3494_re = _RAND_6598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6599 = {1{`RANDOM}};
  _T_3494_im = _RAND_6599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6600 = {1{`RANDOM}};
  _T_3495_re = _RAND_6600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6601 = {1{`RANDOM}};
  _T_3495_im = _RAND_6601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6602 = {1{`RANDOM}};
  _T_3496_re = _RAND_6602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6603 = {1{`RANDOM}};
  _T_3496_im = _RAND_6603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6604 = {1{`RANDOM}};
  _T_3497_re = _RAND_6604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6605 = {1{`RANDOM}};
  _T_3497_im = _RAND_6605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6606 = {1{`RANDOM}};
  _T_3498_re = _RAND_6606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6607 = {1{`RANDOM}};
  _T_3498_im = _RAND_6607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6608 = {1{`RANDOM}};
  _T_3499_re = _RAND_6608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6609 = {1{`RANDOM}};
  _T_3499_im = _RAND_6609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6610 = {1{`RANDOM}};
  _T_3500_re = _RAND_6610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6611 = {1{`RANDOM}};
  _T_3500_im = _RAND_6611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6612 = {1{`RANDOM}};
  _T_3501_re = _RAND_6612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6613 = {1{`RANDOM}};
  _T_3501_im = _RAND_6613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6614 = {1{`RANDOM}};
  _T_3502_re = _RAND_6614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6615 = {1{`RANDOM}};
  _T_3502_im = _RAND_6615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6616 = {1{`RANDOM}};
  _T_3503_re = _RAND_6616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6617 = {1{`RANDOM}};
  _T_3503_im = _RAND_6617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6618 = {1{`RANDOM}};
  _T_3504_re = _RAND_6618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6619 = {1{`RANDOM}};
  _T_3504_im = _RAND_6619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6620 = {1{`RANDOM}};
  _T_3505_re = _RAND_6620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6621 = {1{`RANDOM}};
  _T_3505_im = _RAND_6621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6622 = {1{`RANDOM}};
  _T_3506_re = _RAND_6622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6623 = {1{`RANDOM}};
  _T_3506_im = _RAND_6623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6624 = {1{`RANDOM}};
  _T_3507_re = _RAND_6624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6625 = {1{`RANDOM}};
  _T_3507_im = _RAND_6625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6626 = {1{`RANDOM}};
  _T_3508_re = _RAND_6626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6627 = {1{`RANDOM}};
  _T_3508_im = _RAND_6627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6628 = {1{`RANDOM}};
  _T_3509_re = _RAND_6628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6629 = {1{`RANDOM}};
  _T_3509_im = _RAND_6629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6630 = {1{`RANDOM}};
  _T_3510_re = _RAND_6630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6631 = {1{`RANDOM}};
  _T_3510_im = _RAND_6631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6632 = {1{`RANDOM}};
  _T_3511_re = _RAND_6632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6633 = {1{`RANDOM}};
  _T_3511_im = _RAND_6633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6634 = {1{`RANDOM}};
  _T_3512_re = _RAND_6634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6635 = {1{`RANDOM}};
  _T_3512_im = _RAND_6635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6636 = {1{`RANDOM}};
  _T_3513_re = _RAND_6636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6637 = {1{`RANDOM}};
  _T_3513_im = _RAND_6637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6638 = {1{`RANDOM}};
  _T_3514_re = _RAND_6638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6639 = {1{`RANDOM}};
  _T_3514_im = _RAND_6639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6640 = {1{`RANDOM}};
  _T_3515_re = _RAND_6640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6641 = {1{`RANDOM}};
  _T_3515_im = _RAND_6641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6642 = {1{`RANDOM}};
  _T_3516_re = _RAND_6642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6643 = {1{`RANDOM}};
  _T_3516_im = _RAND_6643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6644 = {1{`RANDOM}};
  _T_3517_re = _RAND_6644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6645 = {1{`RANDOM}};
  _T_3517_im = _RAND_6645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6646 = {1{`RANDOM}};
  _T_3518_re = _RAND_6646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6647 = {1{`RANDOM}};
  _T_3518_im = _RAND_6647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6648 = {1{`RANDOM}};
  _T_3519_re = _RAND_6648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6649 = {1{`RANDOM}};
  _T_3519_im = _RAND_6649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6650 = {1{`RANDOM}};
  _T_3520_re = _RAND_6650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6651 = {1{`RANDOM}};
  _T_3520_im = _RAND_6651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6652 = {1{`RANDOM}};
  _T_3521_re = _RAND_6652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6653 = {1{`RANDOM}};
  _T_3521_im = _RAND_6653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6654 = {1{`RANDOM}};
  _T_3522_re = _RAND_6654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6655 = {1{`RANDOM}};
  _T_3522_im = _RAND_6655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6656 = {1{`RANDOM}};
  _T_3523_re = _RAND_6656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6657 = {1{`RANDOM}};
  _T_3523_im = _RAND_6657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6658 = {1{`RANDOM}};
  _T_3524_re = _RAND_6658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6659 = {1{`RANDOM}};
  _T_3524_im = _RAND_6659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6660 = {1{`RANDOM}};
  _T_3525_re = _RAND_6660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6661 = {1{`RANDOM}};
  _T_3525_im = _RAND_6661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6662 = {1{`RANDOM}};
  _T_3526_re = _RAND_6662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6663 = {1{`RANDOM}};
  _T_3526_im = _RAND_6663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6664 = {1{`RANDOM}};
  _T_3527_re = _RAND_6664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6665 = {1{`RANDOM}};
  _T_3527_im = _RAND_6665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6666 = {1{`RANDOM}};
  _T_3528_re = _RAND_6666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6667 = {1{`RANDOM}};
  _T_3528_im = _RAND_6667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6668 = {1{`RANDOM}};
  _T_3529_re = _RAND_6668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6669 = {1{`RANDOM}};
  _T_3529_im = _RAND_6669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6670 = {1{`RANDOM}};
  _T_3530_re = _RAND_6670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6671 = {1{`RANDOM}};
  _T_3530_im = _RAND_6671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6672 = {1{`RANDOM}};
  _T_3531_re = _RAND_6672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6673 = {1{`RANDOM}};
  _T_3531_im = _RAND_6673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6674 = {1{`RANDOM}};
  _T_3532_re = _RAND_6674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6675 = {1{`RANDOM}};
  _T_3532_im = _RAND_6675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6676 = {1{`RANDOM}};
  _T_3533_re = _RAND_6676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6677 = {1{`RANDOM}};
  _T_3533_im = _RAND_6677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6678 = {1{`RANDOM}};
  _T_3534_re = _RAND_6678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6679 = {1{`RANDOM}};
  _T_3534_im = _RAND_6679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6680 = {1{`RANDOM}};
  _T_3535_re = _RAND_6680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6681 = {1{`RANDOM}};
  _T_3535_im = _RAND_6681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6682 = {1{`RANDOM}};
  _T_3536_re = _RAND_6682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6683 = {1{`RANDOM}};
  _T_3536_im = _RAND_6683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6684 = {1{`RANDOM}};
  _T_3537_re = _RAND_6684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6685 = {1{`RANDOM}};
  _T_3537_im = _RAND_6685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6686 = {1{`RANDOM}};
  _T_3538_re = _RAND_6686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6687 = {1{`RANDOM}};
  _T_3538_im = _RAND_6687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6688 = {1{`RANDOM}};
  _T_3539_re = _RAND_6688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6689 = {1{`RANDOM}};
  _T_3539_im = _RAND_6689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6690 = {1{`RANDOM}};
  _T_3540_re = _RAND_6690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6691 = {1{`RANDOM}};
  _T_3540_im = _RAND_6691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6692 = {1{`RANDOM}};
  _T_3541_re = _RAND_6692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6693 = {1{`RANDOM}};
  _T_3541_im = _RAND_6693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6694 = {1{`RANDOM}};
  _T_3542_re = _RAND_6694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6695 = {1{`RANDOM}};
  _T_3542_im = _RAND_6695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6696 = {1{`RANDOM}};
  _T_3543_re = _RAND_6696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6697 = {1{`RANDOM}};
  _T_3543_im = _RAND_6697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6698 = {1{`RANDOM}};
  _T_3544_re = _RAND_6698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6699 = {1{`RANDOM}};
  _T_3544_im = _RAND_6699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6700 = {1{`RANDOM}};
  _T_3545_re = _RAND_6700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6701 = {1{`RANDOM}};
  _T_3545_im = _RAND_6701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6702 = {1{`RANDOM}};
  _T_3546_re = _RAND_6702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6703 = {1{`RANDOM}};
  _T_3546_im = _RAND_6703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6704 = {1{`RANDOM}};
  _T_3547_re = _RAND_6704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6705 = {1{`RANDOM}};
  _T_3547_im = _RAND_6705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6706 = {1{`RANDOM}};
  _T_3548_re = _RAND_6706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6707 = {1{`RANDOM}};
  _T_3548_im = _RAND_6707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6708 = {1{`RANDOM}};
  _T_3549_re = _RAND_6708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6709 = {1{`RANDOM}};
  _T_3549_im = _RAND_6709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6710 = {1{`RANDOM}};
  _T_3550_re = _RAND_6710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6711 = {1{`RANDOM}};
  _T_3550_im = _RAND_6711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6712 = {1{`RANDOM}};
  _T_3551_re = _RAND_6712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6713 = {1{`RANDOM}};
  _T_3551_im = _RAND_6713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6714 = {1{`RANDOM}};
  _T_3552_re = _RAND_6714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6715 = {1{`RANDOM}};
  _T_3552_im = _RAND_6715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6716 = {1{`RANDOM}};
  _T_3553_re = _RAND_6716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6717 = {1{`RANDOM}};
  _T_3553_im = _RAND_6717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6718 = {1{`RANDOM}};
  _T_3554_re = _RAND_6718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6719 = {1{`RANDOM}};
  _T_3554_im = _RAND_6719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6720 = {1{`RANDOM}};
  _T_3555_re = _RAND_6720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6721 = {1{`RANDOM}};
  _T_3555_im = _RAND_6721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6722 = {1{`RANDOM}};
  _T_3556_re = _RAND_6722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6723 = {1{`RANDOM}};
  _T_3556_im = _RAND_6723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6724 = {1{`RANDOM}};
  _T_3557_re = _RAND_6724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6725 = {1{`RANDOM}};
  _T_3557_im = _RAND_6725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6726 = {1{`RANDOM}};
  _T_3558_re = _RAND_6726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6727 = {1{`RANDOM}};
  _T_3558_im = _RAND_6727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6728 = {1{`RANDOM}};
  _T_3559_re = _RAND_6728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6729 = {1{`RANDOM}};
  _T_3559_im = _RAND_6729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6730 = {1{`RANDOM}};
  _T_3560_re = _RAND_6730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6731 = {1{`RANDOM}};
  _T_3560_im = _RAND_6731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6732 = {1{`RANDOM}};
  _T_3561_re = _RAND_6732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6733 = {1{`RANDOM}};
  _T_3561_im = _RAND_6733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6734 = {1{`RANDOM}};
  _T_3562_re = _RAND_6734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6735 = {1{`RANDOM}};
  _T_3562_im = _RAND_6735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6736 = {1{`RANDOM}};
  _T_3563_re = _RAND_6736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6737 = {1{`RANDOM}};
  _T_3563_im = _RAND_6737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6738 = {1{`RANDOM}};
  _T_3564_re = _RAND_6738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6739 = {1{`RANDOM}};
  _T_3564_im = _RAND_6739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6740 = {1{`RANDOM}};
  _T_3565_re = _RAND_6740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6741 = {1{`RANDOM}};
  _T_3565_im = _RAND_6741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6742 = {1{`RANDOM}};
  _T_3566_re = _RAND_6742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6743 = {1{`RANDOM}};
  _T_3566_im = _RAND_6743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6744 = {1{`RANDOM}};
  _T_3567_re = _RAND_6744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6745 = {1{`RANDOM}};
  _T_3567_im = _RAND_6745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6746 = {1{`RANDOM}};
  _T_3568_re = _RAND_6746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6747 = {1{`RANDOM}};
  _T_3568_im = _RAND_6747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6748 = {1{`RANDOM}};
  _T_3569_re = _RAND_6748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6749 = {1{`RANDOM}};
  _T_3569_im = _RAND_6749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6750 = {1{`RANDOM}};
  _T_3570_re = _RAND_6750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6751 = {1{`RANDOM}};
  _T_3570_im = _RAND_6751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6752 = {1{`RANDOM}};
  _T_3571_re = _RAND_6752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6753 = {1{`RANDOM}};
  _T_3571_im = _RAND_6753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6754 = {1{`RANDOM}};
  _T_3572_re = _RAND_6754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6755 = {1{`RANDOM}};
  _T_3572_im = _RAND_6755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6756 = {1{`RANDOM}};
  _T_3573_re = _RAND_6756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6757 = {1{`RANDOM}};
  _T_3573_im = _RAND_6757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6758 = {1{`RANDOM}};
  _T_3574_re = _RAND_6758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6759 = {1{`RANDOM}};
  _T_3574_im = _RAND_6759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6760 = {1{`RANDOM}};
  _T_3575_re = _RAND_6760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6761 = {1{`RANDOM}};
  _T_3575_im = _RAND_6761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6762 = {1{`RANDOM}};
  _T_3576_re = _RAND_6762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6763 = {1{`RANDOM}};
  _T_3576_im = _RAND_6763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6764 = {1{`RANDOM}};
  _T_3577_re = _RAND_6764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6765 = {1{`RANDOM}};
  _T_3577_im = _RAND_6765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6766 = {1{`RANDOM}};
  _T_3578_re = _RAND_6766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6767 = {1{`RANDOM}};
  _T_3578_im = _RAND_6767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6768 = {1{`RANDOM}};
  _T_3579_re = _RAND_6768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6769 = {1{`RANDOM}};
  _T_3579_im = _RAND_6769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6770 = {1{`RANDOM}};
  _T_3580_re = _RAND_6770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6771 = {1{`RANDOM}};
  _T_3580_im = _RAND_6771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6772 = {1{`RANDOM}};
  _T_3581_re = _RAND_6772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6773 = {1{`RANDOM}};
  _T_3581_im = _RAND_6773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6774 = {1{`RANDOM}};
  _T_3582_re = _RAND_6774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6775 = {1{`RANDOM}};
  _T_3582_im = _RAND_6775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6776 = {1{`RANDOM}};
  _T_3583_re = _RAND_6776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6777 = {1{`RANDOM}};
  _T_3583_im = _RAND_6777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6778 = {1{`RANDOM}};
  _T_3584_re = _RAND_6778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6779 = {1{`RANDOM}};
  _T_3584_im = _RAND_6779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6780 = {1{`RANDOM}};
  _T_3585_re = _RAND_6780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6781 = {1{`RANDOM}};
  _T_3585_im = _RAND_6781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6782 = {1{`RANDOM}};
  _T_3586_re = _RAND_6782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6783 = {1{`RANDOM}};
  _T_3586_im = _RAND_6783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6784 = {1{`RANDOM}};
  _T_3587_re = _RAND_6784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6785 = {1{`RANDOM}};
  _T_3587_im = _RAND_6785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6786 = {1{`RANDOM}};
  _T_3588_re = _RAND_6786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6787 = {1{`RANDOM}};
  _T_3588_im = _RAND_6787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6788 = {1{`RANDOM}};
  _T_3589_re = _RAND_6788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6789 = {1{`RANDOM}};
  _T_3589_im = _RAND_6789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6790 = {1{`RANDOM}};
  _T_3590_re = _RAND_6790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6791 = {1{`RANDOM}};
  _T_3590_im = _RAND_6791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6792 = {1{`RANDOM}};
  _T_3591_re = _RAND_6792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6793 = {1{`RANDOM}};
  _T_3591_im = _RAND_6793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6794 = {1{`RANDOM}};
  _T_3592_re = _RAND_6794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6795 = {1{`RANDOM}};
  _T_3592_im = _RAND_6795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6796 = {1{`RANDOM}};
  _T_3593_re = _RAND_6796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6797 = {1{`RANDOM}};
  _T_3593_im = _RAND_6797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6798 = {1{`RANDOM}};
  _T_3594_re = _RAND_6798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6799 = {1{`RANDOM}};
  _T_3594_im = _RAND_6799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6800 = {1{`RANDOM}};
  _T_3595_re = _RAND_6800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6801 = {1{`RANDOM}};
  _T_3595_im = _RAND_6801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6802 = {1{`RANDOM}};
  _T_3596_re = _RAND_6802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6803 = {1{`RANDOM}};
  _T_3596_im = _RAND_6803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6804 = {1{`RANDOM}};
  _T_3597_re = _RAND_6804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6805 = {1{`RANDOM}};
  _T_3597_im = _RAND_6805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6806 = {1{`RANDOM}};
  _T_3598_re = _RAND_6806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6807 = {1{`RANDOM}};
  _T_3598_im = _RAND_6807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6808 = {1{`RANDOM}};
  _T_3599_re = _RAND_6808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6809 = {1{`RANDOM}};
  _T_3599_im = _RAND_6809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6810 = {1{`RANDOM}};
  _T_3600_re = _RAND_6810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6811 = {1{`RANDOM}};
  _T_3600_im = _RAND_6811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6812 = {1{`RANDOM}};
  _T_3601_re = _RAND_6812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6813 = {1{`RANDOM}};
  _T_3601_im = _RAND_6813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6814 = {1{`RANDOM}};
  _T_3602_re = _RAND_6814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6815 = {1{`RANDOM}};
  _T_3602_im = _RAND_6815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6816 = {1{`RANDOM}};
  _T_3603_re = _RAND_6816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6817 = {1{`RANDOM}};
  _T_3603_im = _RAND_6817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6818 = {1{`RANDOM}};
  _T_3604_re = _RAND_6818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6819 = {1{`RANDOM}};
  _T_3604_im = _RAND_6819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6820 = {1{`RANDOM}};
  _T_3605_re = _RAND_6820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6821 = {1{`RANDOM}};
  _T_3605_im = _RAND_6821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6822 = {1{`RANDOM}};
  _T_3606_re = _RAND_6822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6823 = {1{`RANDOM}};
  _T_3606_im = _RAND_6823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6824 = {1{`RANDOM}};
  _T_3607_re = _RAND_6824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6825 = {1{`RANDOM}};
  _T_3607_im = _RAND_6825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6826 = {1{`RANDOM}};
  _T_3608_re = _RAND_6826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6827 = {1{`RANDOM}};
  _T_3608_im = _RAND_6827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6828 = {1{`RANDOM}};
  _T_3609_re = _RAND_6828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6829 = {1{`RANDOM}};
  _T_3609_im = _RAND_6829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6830 = {1{`RANDOM}};
  _T_3610_re = _RAND_6830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6831 = {1{`RANDOM}};
  _T_3610_im = _RAND_6831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6832 = {1{`RANDOM}};
  _T_3611_re = _RAND_6832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6833 = {1{`RANDOM}};
  _T_3611_im = _RAND_6833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6834 = {1{`RANDOM}};
  _T_3612_re = _RAND_6834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6835 = {1{`RANDOM}};
  _T_3612_im = _RAND_6835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6836 = {1{`RANDOM}};
  _T_3613_re = _RAND_6836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6837 = {1{`RANDOM}};
  _T_3613_im = _RAND_6837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6838 = {1{`RANDOM}};
  _T_3614_re = _RAND_6838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6839 = {1{`RANDOM}};
  _T_3614_im = _RAND_6839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6840 = {1{`RANDOM}};
  _T_3615_re = _RAND_6840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6841 = {1{`RANDOM}};
  _T_3615_im = _RAND_6841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6842 = {1{`RANDOM}};
  _T_3616_re = _RAND_6842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6843 = {1{`RANDOM}};
  _T_3616_im = _RAND_6843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6844 = {1{`RANDOM}};
  _T_3617_re = _RAND_6844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6845 = {1{`RANDOM}};
  _T_3617_im = _RAND_6845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6846 = {1{`RANDOM}};
  _T_3618_re = _RAND_6846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6847 = {1{`RANDOM}};
  _T_3618_im = _RAND_6847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6848 = {1{`RANDOM}};
  _T_3619_re = _RAND_6848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6849 = {1{`RANDOM}};
  _T_3619_im = _RAND_6849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6850 = {1{`RANDOM}};
  _T_3620_re = _RAND_6850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6851 = {1{`RANDOM}};
  _T_3620_im = _RAND_6851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6852 = {1{`RANDOM}};
  _T_3621_re = _RAND_6852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6853 = {1{`RANDOM}};
  _T_3621_im = _RAND_6853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6854 = {1{`RANDOM}};
  _T_3622_re = _RAND_6854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6855 = {1{`RANDOM}};
  _T_3622_im = _RAND_6855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6856 = {1{`RANDOM}};
  _T_3623_re = _RAND_6856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6857 = {1{`RANDOM}};
  _T_3623_im = _RAND_6857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6858 = {1{`RANDOM}};
  _T_3624_re = _RAND_6858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6859 = {1{`RANDOM}};
  _T_3624_im = _RAND_6859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6860 = {1{`RANDOM}};
  _T_3625_re = _RAND_6860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6861 = {1{`RANDOM}};
  _T_3625_im = _RAND_6861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6862 = {1{`RANDOM}};
  _T_3626_re = _RAND_6862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6863 = {1{`RANDOM}};
  _T_3626_im = _RAND_6863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6864 = {1{`RANDOM}};
  _T_3627_re = _RAND_6864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6865 = {1{`RANDOM}};
  _T_3627_im = _RAND_6865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6866 = {1{`RANDOM}};
  _T_3628_re = _RAND_6866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6867 = {1{`RANDOM}};
  _T_3628_im = _RAND_6867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6868 = {1{`RANDOM}};
  _T_3629_re = _RAND_6868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6869 = {1{`RANDOM}};
  _T_3629_im = _RAND_6869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6870 = {1{`RANDOM}};
  _T_3630_re = _RAND_6870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6871 = {1{`RANDOM}};
  _T_3630_im = _RAND_6871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6872 = {1{`RANDOM}};
  _T_3631_re = _RAND_6872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6873 = {1{`RANDOM}};
  _T_3631_im = _RAND_6873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6874 = {1{`RANDOM}};
  _T_3632_re = _RAND_6874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6875 = {1{`RANDOM}};
  _T_3632_im = _RAND_6875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6876 = {1{`RANDOM}};
  _T_3633_re = _RAND_6876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6877 = {1{`RANDOM}};
  _T_3633_im = _RAND_6877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6878 = {1{`RANDOM}};
  _T_3634_re = _RAND_6878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6879 = {1{`RANDOM}};
  _T_3634_im = _RAND_6879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6880 = {1{`RANDOM}};
  _T_3635_re = _RAND_6880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6881 = {1{`RANDOM}};
  _T_3635_im = _RAND_6881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6882 = {1{`RANDOM}};
  _T_3636_re = _RAND_6882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6883 = {1{`RANDOM}};
  _T_3636_im = _RAND_6883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6884 = {1{`RANDOM}};
  _T_3637_re = _RAND_6884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6885 = {1{`RANDOM}};
  _T_3637_im = _RAND_6885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6886 = {1{`RANDOM}};
  _T_3638_re = _RAND_6886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6887 = {1{`RANDOM}};
  _T_3638_im = _RAND_6887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6888 = {1{`RANDOM}};
  _T_3639_re = _RAND_6888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6889 = {1{`RANDOM}};
  _T_3639_im = _RAND_6889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6890 = {1{`RANDOM}};
  _T_3640_re = _RAND_6890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6891 = {1{`RANDOM}};
  _T_3640_im = _RAND_6891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6892 = {1{`RANDOM}};
  _T_3641_re = _RAND_6892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6893 = {1{`RANDOM}};
  _T_3641_im = _RAND_6893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6894 = {1{`RANDOM}};
  _T_3642_re = _RAND_6894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6895 = {1{`RANDOM}};
  _T_3642_im = _RAND_6895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6896 = {1{`RANDOM}};
  _T_3643_re = _RAND_6896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6897 = {1{`RANDOM}};
  _T_3643_im = _RAND_6897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6898 = {1{`RANDOM}};
  _T_3644_re = _RAND_6898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6899 = {1{`RANDOM}};
  _T_3644_im = _RAND_6899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6900 = {1{`RANDOM}};
  _T_3645_re = _RAND_6900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6901 = {1{`RANDOM}};
  _T_3645_im = _RAND_6901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6902 = {1{`RANDOM}};
  _T_3646_re = _RAND_6902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6903 = {1{`RANDOM}};
  _T_3646_im = _RAND_6903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6904 = {1{`RANDOM}};
  _T_3647_re = _RAND_6904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6905 = {1{`RANDOM}};
  _T_3647_im = _RAND_6905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6906 = {1{`RANDOM}};
  _T_3648_re = _RAND_6906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6907 = {1{`RANDOM}};
  _T_3648_im = _RAND_6907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6908 = {1{`RANDOM}};
  _T_3649_re = _RAND_6908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6909 = {1{`RANDOM}};
  _T_3649_im = _RAND_6909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6910 = {1{`RANDOM}};
  _T_3650_re = _RAND_6910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6911 = {1{`RANDOM}};
  _T_3650_im = _RAND_6911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6912 = {1{`RANDOM}};
  _T_3651_re = _RAND_6912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6913 = {1{`RANDOM}};
  _T_3651_im = _RAND_6913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6914 = {1{`RANDOM}};
  _T_3652_re = _RAND_6914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6915 = {1{`RANDOM}};
  _T_3652_im = _RAND_6915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6916 = {1{`RANDOM}};
  _T_3653_re = _RAND_6916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6917 = {1{`RANDOM}};
  _T_3653_im = _RAND_6917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6918 = {1{`RANDOM}};
  _T_3654_re = _RAND_6918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6919 = {1{`RANDOM}};
  _T_3654_im = _RAND_6919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6920 = {1{`RANDOM}};
  _T_3655_re = _RAND_6920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6921 = {1{`RANDOM}};
  _T_3655_im = _RAND_6921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6922 = {1{`RANDOM}};
  _T_3656_re = _RAND_6922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6923 = {1{`RANDOM}};
  _T_3656_im = _RAND_6923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6924 = {1{`RANDOM}};
  _T_3657_re = _RAND_6924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6925 = {1{`RANDOM}};
  _T_3657_im = _RAND_6925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6926 = {1{`RANDOM}};
  _T_3658_re = _RAND_6926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6927 = {1{`RANDOM}};
  _T_3658_im = _RAND_6927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6928 = {1{`RANDOM}};
  _T_3659_re = _RAND_6928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6929 = {1{`RANDOM}};
  _T_3659_im = _RAND_6929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6930 = {1{`RANDOM}};
  _T_3660_re = _RAND_6930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6931 = {1{`RANDOM}};
  _T_3660_im = _RAND_6931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6932 = {1{`RANDOM}};
  _T_3661_re = _RAND_6932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6933 = {1{`RANDOM}};
  _T_3661_im = _RAND_6933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6934 = {1{`RANDOM}};
  _T_3662_re = _RAND_6934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6935 = {1{`RANDOM}};
  _T_3662_im = _RAND_6935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6936 = {1{`RANDOM}};
  _T_3663_re = _RAND_6936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6937 = {1{`RANDOM}};
  _T_3663_im = _RAND_6937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6938 = {1{`RANDOM}};
  _T_3664_re = _RAND_6938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6939 = {1{`RANDOM}};
  _T_3664_im = _RAND_6939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6940 = {1{`RANDOM}};
  _T_3665_re = _RAND_6940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6941 = {1{`RANDOM}};
  _T_3665_im = _RAND_6941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6942 = {1{`RANDOM}};
  _T_3666_re = _RAND_6942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6943 = {1{`RANDOM}};
  _T_3666_im = _RAND_6943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6944 = {1{`RANDOM}};
  _T_3667_re = _RAND_6944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6945 = {1{`RANDOM}};
  _T_3667_im = _RAND_6945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6946 = {1{`RANDOM}};
  _T_3668_re = _RAND_6946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6947 = {1{`RANDOM}};
  _T_3668_im = _RAND_6947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6948 = {1{`RANDOM}};
  _T_3669_re = _RAND_6948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6949 = {1{`RANDOM}};
  _T_3669_im = _RAND_6949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6950 = {1{`RANDOM}};
  _T_3670_re = _RAND_6950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6951 = {1{`RANDOM}};
  _T_3670_im = _RAND_6951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6952 = {1{`RANDOM}};
  _T_3671_re = _RAND_6952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6953 = {1{`RANDOM}};
  _T_3671_im = _RAND_6953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6954 = {1{`RANDOM}};
  _T_3672_re = _RAND_6954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6955 = {1{`RANDOM}};
  _T_3672_im = _RAND_6955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6956 = {1{`RANDOM}};
  _T_3673_re = _RAND_6956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6957 = {1{`RANDOM}};
  _T_3673_im = _RAND_6957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6958 = {1{`RANDOM}};
  _T_3674_re = _RAND_6958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6959 = {1{`RANDOM}};
  _T_3674_im = _RAND_6959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6960 = {1{`RANDOM}};
  _T_3675_re = _RAND_6960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6961 = {1{`RANDOM}};
  _T_3675_im = _RAND_6961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6962 = {1{`RANDOM}};
  _T_3676_re = _RAND_6962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6963 = {1{`RANDOM}};
  _T_3676_im = _RAND_6963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6964 = {1{`RANDOM}};
  _T_3677_re = _RAND_6964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6965 = {1{`RANDOM}};
  _T_3677_im = _RAND_6965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6966 = {1{`RANDOM}};
  _T_3678_re = _RAND_6966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6967 = {1{`RANDOM}};
  _T_3678_im = _RAND_6967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6968 = {1{`RANDOM}};
  _T_3679_re = _RAND_6968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6969 = {1{`RANDOM}};
  _T_3679_im = _RAND_6969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6970 = {1{`RANDOM}};
  _T_3680_re = _RAND_6970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6971 = {1{`RANDOM}};
  _T_3680_im = _RAND_6971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6972 = {1{`RANDOM}};
  _T_3681_re = _RAND_6972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6973 = {1{`RANDOM}};
  _T_3681_im = _RAND_6973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6974 = {1{`RANDOM}};
  _T_3682_re = _RAND_6974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6975 = {1{`RANDOM}};
  _T_3682_im = _RAND_6975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6976 = {1{`RANDOM}};
  _T_3683_re = _RAND_6976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6977 = {1{`RANDOM}};
  _T_3683_im = _RAND_6977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6978 = {1{`RANDOM}};
  _T_3684_re = _RAND_6978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6979 = {1{`RANDOM}};
  _T_3684_im = _RAND_6979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6980 = {1{`RANDOM}};
  _T_3685_re = _RAND_6980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6981 = {1{`RANDOM}};
  _T_3685_im = _RAND_6981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6982 = {1{`RANDOM}};
  _T_3686_re = _RAND_6982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6983 = {1{`RANDOM}};
  _T_3686_im = _RAND_6983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6984 = {1{`RANDOM}};
  _T_3687_re = _RAND_6984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6985 = {1{`RANDOM}};
  _T_3687_im = _RAND_6985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6986 = {1{`RANDOM}};
  _T_3688_re = _RAND_6986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6987 = {1{`RANDOM}};
  _T_3688_im = _RAND_6987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6988 = {1{`RANDOM}};
  _T_3689_re = _RAND_6988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6989 = {1{`RANDOM}};
  _T_3689_im = _RAND_6989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6990 = {1{`RANDOM}};
  _T_3690_re = _RAND_6990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6991 = {1{`RANDOM}};
  _T_3690_im = _RAND_6991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6992 = {1{`RANDOM}};
  _T_3691_re = _RAND_6992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6993 = {1{`RANDOM}};
  _T_3691_im = _RAND_6993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6994 = {1{`RANDOM}};
  _T_3692_re = _RAND_6994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6995 = {1{`RANDOM}};
  _T_3692_im = _RAND_6995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6996 = {1{`RANDOM}};
  _T_3693_re = _RAND_6996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6997 = {1{`RANDOM}};
  _T_3693_im = _RAND_6997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6998 = {1{`RANDOM}};
  _T_3694_re = _RAND_6998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6999 = {1{`RANDOM}};
  _T_3694_im = _RAND_6999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7000 = {1{`RANDOM}};
  _T_3695_re = _RAND_7000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7001 = {1{`RANDOM}};
  _T_3695_im = _RAND_7001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7002 = {1{`RANDOM}};
  _T_3696_re = _RAND_7002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7003 = {1{`RANDOM}};
  _T_3696_im = _RAND_7003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7004 = {1{`RANDOM}};
  _T_3697_re = _RAND_7004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7005 = {1{`RANDOM}};
  _T_3697_im = _RAND_7005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7006 = {1{`RANDOM}};
  _T_3698_re = _RAND_7006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7007 = {1{`RANDOM}};
  _T_3698_im = _RAND_7007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7008 = {1{`RANDOM}};
  _T_3699_re = _RAND_7008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7009 = {1{`RANDOM}};
  _T_3699_im = _RAND_7009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7010 = {1{`RANDOM}};
  _T_3700_re = _RAND_7010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7011 = {1{`RANDOM}};
  _T_3700_im = _RAND_7011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7012 = {1{`RANDOM}};
  _T_3701_re = _RAND_7012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7013 = {1{`RANDOM}};
  _T_3701_im = _RAND_7013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7014 = {1{`RANDOM}};
  _T_3702_re = _RAND_7014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7015 = {1{`RANDOM}};
  _T_3702_im = _RAND_7015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7016 = {1{`RANDOM}};
  _T_3703_re = _RAND_7016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7017 = {1{`RANDOM}};
  _T_3703_im = _RAND_7017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7018 = {1{`RANDOM}};
  _T_3704_re = _RAND_7018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7019 = {1{`RANDOM}};
  _T_3704_im = _RAND_7019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7020 = {1{`RANDOM}};
  _T_3705_re = _RAND_7020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7021 = {1{`RANDOM}};
  _T_3705_im = _RAND_7021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7022 = {1{`RANDOM}};
  _T_3706_re = _RAND_7022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7023 = {1{`RANDOM}};
  _T_3706_im = _RAND_7023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7024 = {1{`RANDOM}};
  _T_3707_re = _RAND_7024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7025 = {1{`RANDOM}};
  _T_3707_im = _RAND_7025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7026 = {1{`RANDOM}};
  _T_3708_re = _RAND_7026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7027 = {1{`RANDOM}};
  _T_3708_im = _RAND_7027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7028 = {1{`RANDOM}};
  _T_3709_re = _RAND_7028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7029 = {1{`RANDOM}};
  _T_3709_im = _RAND_7029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7030 = {1{`RANDOM}};
  _T_3710_re = _RAND_7030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7031 = {1{`RANDOM}};
  _T_3710_im = _RAND_7031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7032 = {1{`RANDOM}};
  _T_3711_re = _RAND_7032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7033 = {1{`RANDOM}};
  _T_3711_im = _RAND_7033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7034 = {1{`RANDOM}};
  _T_3712_re = _RAND_7034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7035 = {1{`RANDOM}};
  _T_3712_im = _RAND_7035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7036 = {1{`RANDOM}};
  _T_3713_re = _RAND_7036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7037 = {1{`RANDOM}};
  _T_3713_im = _RAND_7037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7038 = {1{`RANDOM}};
  _T_3714_re = _RAND_7038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7039 = {1{`RANDOM}};
  _T_3714_im = _RAND_7039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7040 = {1{`RANDOM}};
  _T_3715_re = _RAND_7040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7041 = {1{`RANDOM}};
  _T_3715_im = _RAND_7041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7042 = {1{`RANDOM}};
  _T_3716_re = _RAND_7042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7043 = {1{`RANDOM}};
  _T_3716_im = _RAND_7043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7044 = {1{`RANDOM}};
  _T_3717_re = _RAND_7044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7045 = {1{`RANDOM}};
  _T_3717_im = _RAND_7045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7046 = {1{`RANDOM}};
  _T_3718_re = _RAND_7046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7047 = {1{`RANDOM}};
  _T_3718_im = _RAND_7047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7048 = {1{`RANDOM}};
  _T_3719_re = _RAND_7048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7049 = {1{`RANDOM}};
  _T_3719_im = _RAND_7049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7050 = {1{`RANDOM}};
  _T_3720_re = _RAND_7050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7051 = {1{`RANDOM}};
  _T_3720_im = _RAND_7051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7052 = {1{`RANDOM}};
  _T_3721_re = _RAND_7052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7053 = {1{`RANDOM}};
  _T_3721_im = _RAND_7053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7054 = {1{`RANDOM}};
  _T_3722_re = _RAND_7054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7055 = {1{`RANDOM}};
  _T_3722_im = _RAND_7055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7056 = {1{`RANDOM}};
  _T_3723_re = _RAND_7056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7057 = {1{`RANDOM}};
  _T_3723_im = _RAND_7057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7058 = {1{`RANDOM}};
  _T_3724_re = _RAND_7058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7059 = {1{`RANDOM}};
  _T_3724_im = _RAND_7059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7060 = {1{`RANDOM}};
  _T_3725_re = _RAND_7060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7061 = {1{`RANDOM}};
  _T_3725_im = _RAND_7061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7062 = {1{`RANDOM}};
  _T_3726_re = _RAND_7062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7063 = {1{`RANDOM}};
  _T_3726_im = _RAND_7063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7064 = {1{`RANDOM}};
  _T_3727_re = _RAND_7064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7065 = {1{`RANDOM}};
  _T_3727_im = _RAND_7065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7066 = {1{`RANDOM}};
  _T_3728_re = _RAND_7066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7067 = {1{`RANDOM}};
  _T_3728_im = _RAND_7067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7068 = {1{`RANDOM}};
  _T_3729_re = _RAND_7068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7069 = {1{`RANDOM}};
  _T_3729_im = _RAND_7069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7070 = {1{`RANDOM}};
  _T_3730_re = _RAND_7070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7071 = {1{`RANDOM}};
  _T_3730_im = _RAND_7071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7072 = {1{`RANDOM}};
  _T_3731_re = _RAND_7072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7073 = {1{`RANDOM}};
  _T_3731_im = _RAND_7073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7074 = {1{`RANDOM}};
  _T_3732_re = _RAND_7074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7075 = {1{`RANDOM}};
  _T_3732_im = _RAND_7075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7076 = {1{`RANDOM}};
  _T_3733_re = _RAND_7076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7077 = {1{`RANDOM}};
  _T_3733_im = _RAND_7077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7078 = {1{`RANDOM}};
  _T_3734_re = _RAND_7078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7079 = {1{`RANDOM}};
  _T_3734_im = _RAND_7079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7080 = {1{`RANDOM}};
  _T_3735_re = _RAND_7080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7081 = {1{`RANDOM}};
  _T_3735_im = _RAND_7081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7082 = {1{`RANDOM}};
  _T_3736_re = _RAND_7082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7083 = {1{`RANDOM}};
  _T_3736_im = _RAND_7083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7084 = {1{`RANDOM}};
  _T_3737_re = _RAND_7084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7085 = {1{`RANDOM}};
  _T_3737_im = _RAND_7085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7086 = {1{`RANDOM}};
  _T_3738_re = _RAND_7086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7087 = {1{`RANDOM}};
  _T_3738_im = _RAND_7087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7088 = {1{`RANDOM}};
  _T_3739_re = _RAND_7088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7089 = {1{`RANDOM}};
  _T_3739_im = _RAND_7089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7090 = {1{`RANDOM}};
  _T_3740_re = _RAND_7090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7091 = {1{`RANDOM}};
  _T_3740_im = _RAND_7091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7092 = {1{`RANDOM}};
  _T_3741_re = _RAND_7092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7093 = {1{`RANDOM}};
  _T_3741_im = _RAND_7093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7094 = {1{`RANDOM}};
  _T_3742_re = _RAND_7094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7095 = {1{`RANDOM}};
  _T_3742_im = _RAND_7095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7096 = {1{`RANDOM}};
  _T_3743_re = _RAND_7096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7097 = {1{`RANDOM}};
  _T_3743_im = _RAND_7097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7098 = {1{`RANDOM}};
  _T_3744_re = _RAND_7098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7099 = {1{`RANDOM}};
  _T_3744_im = _RAND_7099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7100 = {1{`RANDOM}};
  _T_3745_re = _RAND_7100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7101 = {1{`RANDOM}};
  _T_3745_im = _RAND_7101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7102 = {1{`RANDOM}};
  _T_3746_re = _RAND_7102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7103 = {1{`RANDOM}};
  _T_3746_im = _RAND_7103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7104 = {1{`RANDOM}};
  _T_3747_re = _RAND_7104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7105 = {1{`RANDOM}};
  _T_3747_im = _RAND_7105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7106 = {1{`RANDOM}};
  _T_3748_re = _RAND_7106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7107 = {1{`RANDOM}};
  _T_3748_im = _RAND_7107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7108 = {1{`RANDOM}};
  _T_3749_re = _RAND_7108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7109 = {1{`RANDOM}};
  _T_3749_im = _RAND_7109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7110 = {1{`RANDOM}};
  _T_3750_re = _RAND_7110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7111 = {1{`RANDOM}};
  _T_3750_im = _RAND_7111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7112 = {1{`RANDOM}};
  _T_3751_re = _RAND_7112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7113 = {1{`RANDOM}};
  _T_3751_im = _RAND_7113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7114 = {1{`RANDOM}};
  _T_3752_re = _RAND_7114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7115 = {1{`RANDOM}};
  _T_3752_im = _RAND_7115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7116 = {1{`RANDOM}};
  _T_3753_re = _RAND_7116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7117 = {1{`RANDOM}};
  _T_3753_im = _RAND_7117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7118 = {1{`RANDOM}};
  _T_3754_re = _RAND_7118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7119 = {1{`RANDOM}};
  _T_3754_im = _RAND_7119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7120 = {1{`RANDOM}};
  _T_3755_re = _RAND_7120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7121 = {1{`RANDOM}};
  _T_3755_im = _RAND_7121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7122 = {1{`RANDOM}};
  _T_3756_re = _RAND_7122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7123 = {1{`RANDOM}};
  _T_3756_im = _RAND_7123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7124 = {1{`RANDOM}};
  _T_3757_re = _RAND_7124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7125 = {1{`RANDOM}};
  _T_3757_im = _RAND_7125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7126 = {1{`RANDOM}};
  _T_3758_re = _RAND_7126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7127 = {1{`RANDOM}};
  _T_3758_im = _RAND_7127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7128 = {1{`RANDOM}};
  _T_3759_re = _RAND_7128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7129 = {1{`RANDOM}};
  _T_3759_im = _RAND_7129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7130 = {1{`RANDOM}};
  _T_3760_re = _RAND_7130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7131 = {1{`RANDOM}};
  _T_3760_im = _RAND_7131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7132 = {1{`RANDOM}};
  _T_3761_re = _RAND_7132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7133 = {1{`RANDOM}};
  _T_3761_im = _RAND_7133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7134 = {1{`RANDOM}};
  _T_3762_re = _RAND_7134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7135 = {1{`RANDOM}};
  _T_3762_im = _RAND_7135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7136 = {1{`RANDOM}};
  _T_3763_re = _RAND_7136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7137 = {1{`RANDOM}};
  _T_3763_im = _RAND_7137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7138 = {1{`RANDOM}};
  _T_3764_re = _RAND_7138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7139 = {1{`RANDOM}};
  _T_3764_im = _RAND_7139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7140 = {1{`RANDOM}};
  _T_3765_re = _RAND_7140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7141 = {1{`RANDOM}};
  _T_3765_im = _RAND_7141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7142 = {1{`RANDOM}};
  _T_3766_re = _RAND_7142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7143 = {1{`RANDOM}};
  _T_3766_im = _RAND_7143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7144 = {1{`RANDOM}};
  _T_3767_re = _RAND_7144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7145 = {1{`RANDOM}};
  _T_3767_im = _RAND_7145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7146 = {1{`RANDOM}};
  _T_3768_re = _RAND_7146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7147 = {1{`RANDOM}};
  _T_3768_im = _RAND_7147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7148 = {1{`RANDOM}};
  _T_3769_re = _RAND_7148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7149 = {1{`RANDOM}};
  _T_3769_im = _RAND_7149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7150 = {1{`RANDOM}};
  _T_3770_re = _RAND_7150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7151 = {1{`RANDOM}};
  _T_3770_im = _RAND_7151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7152 = {1{`RANDOM}};
  _T_3771_re = _RAND_7152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7153 = {1{`RANDOM}};
  _T_3771_im = _RAND_7153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7154 = {1{`RANDOM}};
  _T_3772_re = _RAND_7154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7155 = {1{`RANDOM}};
  _T_3772_im = _RAND_7155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7156 = {1{`RANDOM}};
  _T_3773_re = _RAND_7156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7157 = {1{`RANDOM}};
  _T_3773_im = _RAND_7157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7158 = {1{`RANDOM}};
  _T_3774_re = _RAND_7158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7159 = {1{`RANDOM}};
  _T_3774_im = _RAND_7159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7160 = {1{`RANDOM}};
  _T_3775_re = _RAND_7160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7161 = {1{`RANDOM}};
  _T_3775_im = _RAND_7161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7162 = {1{`RANDOM}};
  _T_3776_re = _RAND_7162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7163 = {1{`RANDOM}};
  _T_3776_im = _RAND_7163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7164 = {1{`RANDOM}};
  _T_3777_re = _RAND_7164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7165 = {1{`RANDOM}};
  _T_3777_im = _RAND_7165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7166 = {1{`RANDOM}};
  _T_3778_re = _RAND_7166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7167 = {1{`RANDOM}};
  _T_3778_im = _RAND_7167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7168 = {1{`RANDOM}};
  _T_3779_re = _RAND_7168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7169 = {1{`RANDOM}};
  _T_3779_im = _RAND_7169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7170 = {1{`RANDOM}};
  _T_3780_re = _RAND_7170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7171 = {1{`RANDOM}};
  _T_3780_im = _RAND_7171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7172 = {1{`RANDOM}};
  _T_3781_re = _RAND_7172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7173 = {1{`RANDOM}};
  _T_3781_im = _RAND_7173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7174 = {1{`RANDOM}};
  _T_3782_re = _RAND_7174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7175 = {1{`RANDOM}};
  _T_3782_im = _RAND_7175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7176 = {1{`RANDOM}};
  _T_3783_re = _RAND_7176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7177 = {1{`RANDOM}};
  _T_3783_im = _RAND_7177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7178 = {1{`RANDOM}};
  _T_3784_re = _RAND_7178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7179 = {1{`RANDOM}};
  _T_3784_im = _RAND_7179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7180 = {1{`RANDOM}};
  _T_3785_re = _RAND_7180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7181 = {1{`RANDOM}};
  _T_3785_im = _RAND_7181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7182 = {1{`RANDOM}};
  _T_3786_re = _RAND_7182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7183 = {1{`RANDOM}};
  _T_3786_im = _RAND_7183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7184 = {1{`RANDOM}};
  _T_3787_re = _RAND_7184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7185 = {1{`RANDOM}};
  _T_3787_im = _RAND_7185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7186 = {1{`RANDOM}};
  _T_3788_re = _RAND_7186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7187 = {1{`RANDOM}};
  _T_3788_im = _RAND_7187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7188 = {1{`RANDOM}};
  _T_3789_re = _RAND_7188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7189 = {1{`RANDOM}};
  _T_3789_im = _RAND_7189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7190 = {1{`RANDOM}};
  _T_3790_re = _RAND_7190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7191 = {1{`RANDOM}};
  _T_3790_im = _RAND_7191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7192 = {1{`RANDOM}};
  _T_3791_re = _RAND_7192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7193 = {1{`RANDOM}};
  _T_3791_im = _RAND_7193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7194 = {1{`RANDOM}};
  _T_3792_re = _RAND_7194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7195 = {1{`RANDOM}};
  _T_3792_im = _RAND_7195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7196 = {1{`RANDOM}};
  _T_3793_re = _RAND_7196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7197 = {1{`RANDOM}};
  _T_3793_im = _RAND_7197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7198 = {1{`RANDOM}};
  _T_3794_re = _RAND_7198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7199 = {1{`RANDOM}};
  _T_3794_im = _RAND_7199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7200 = {1{`RANDOM}};
  _T_3795_re = _RAND_7200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7201 = {1{`RANDOM}};
  _T_3795_im = _RAND_7201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7202 = {1{`RANDOM}};
  _T_3796_re = _RAND_7202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7203 = {1{`RANDOM}};
  _T_3796_im = _RAND_7203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7204 = {1{`RANDOM}};
  _T_3797_re = _RAND_7204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7205 = {1{`RANDOM}};
  _T_3797_im = _RAND_7205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7206 = {1{`RANDOM}};
  _T_3798_re = _RAND_7206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7207 = {1{`RANDOM}};
  _T_3798_im = _RAND_7207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7208 = {1{`RANDOM}};
  _T_3799_re = _RAND_7208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7209 = {1{`RANDOM}};
  _T_3799_im = _RAND_7209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7210 = {1{`RANDOM}};
  _T_3800_re = _RAND_7210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7211 = {1{`RANDOM}};
  _T_3800_im = _RAND_7211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7212 = {1{`RANDOM}};
  _T_3801_re = _RAND_7212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7213 = {1{`RANDOM}};
  _T_3801_im = _RAND_7213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7214 = {1{`RANDOM}};
  _T_3802_re = _RAND_7214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7215 = {1{`RANDOM}};
  _T_3802_im = _RAND_7215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7216 = {1{`RANDOM}};
  _T_3803_re = _RAND_7216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7217 = {1{`RANDOM}};
  _T_3803_im = _RAND_7217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7218 = {1{`RANDOM}};
  _T_3804_re = _RAND_7218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7219 = {1{`RANDOM}};
  _T_3804_im = _RAND_7219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7220 = {1{`RANDOM}};
  _T_3805_re = _RAND_7220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7221 = {1{`RANDOM}};
  _T_3805_im = _RAND_7221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7222 = {1{`RANDOM}};
  _T_3806_re = _RAND_7222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7223 = {1{`RANDOM}};
  _T_3806_im = _RAND_7223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7224 = {1{`RANDOM}};
  _T_3807_re = _RAND_7224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7225 = {1{`RANDOM}};
  _T_3807_im = _RAND_7225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7226 = {1{`RANDOM}};
  _T_3808_re = _RAND_7226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7227 = {1{`RANDOM}};
  _T_3808_im = _RAND_7227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7228 = {1{`RANDOM}};
  _T_3809_re = _RAND_7228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7229 = {1{`RANDOM}};
  _T_3809_im = _RAND_7229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7230 = {1{`RANDOM}};
  _T_3810_re = _RAND_7230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7231 = {1{`RANDOM}};
  _T_3810_im = _RAND_7231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7232 = {1{`RANDOM}};
  _T_3811_re = _RAND_7232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7233 = {1{`RANDOM}};
  _T_3811_im = _RAND_7233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7234 = {1{`RANDOM}};
  _T_3812_re = _RAND_7234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7235 = {1{`RANDOM}};
  _T_3812_im = _RAND_7235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7236 = {1{`RANDOM}};
  _T_3813_re = _RAND_7236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7237 = {1{`RANDOM}};
  _T_3813_im = _RAND_7237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7238 = {1{`RANDOM}};
  _T_3814_re = _RAND_7238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7239 = {1{`RANDOM}};
  _T_3814_im = _RAND_7239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7240 = {1{`RANDOM}};
  _T_3815_re = _RAND_7240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7241 = {1{`RANDOM}};
  _T_3815_im = _RAND_7241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7242 = {1{`RANDOM}};
  _T_3816_re = _RAND_7242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7243 = {1{`RANDOM}};
  _T_3816_im = _RAND_7243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7244 = {1{`RANDOM}};
  _T_3817_re = _RAND_7244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7245 = {1{`RANDOM}};
  _T_3817_im = _RAND_7245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7246 = {1{`RANDOM}};
  _T_3818_re = _RAND_7246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7247 = {1{`RANDOM}};
  _T_3818_im = _RAND_7247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7248 = {1{`RANDOM}};
  _T_3819_re = _RAND_7248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7249 = {1{`RANDOM}};
  _T_3819_im = _RAND_7249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7250 = {1{`RANDOM}};
  _T_3820_re = _RAND_7250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7251 = {1{`RANDOM}};
  _T_3820_im = _RAND_7251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7252 = {1{`RANDOM}};
  _T_3821_re = _RAND_7252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7253 = {1{`RANDOM}};
  _T_3821_im = _RAND_7253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7254 = {1{`RANDOM}};
  _T_3822_re = _RAND_7254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7255 = {1{`RANDOM}};
  _T_3822_im = _RAND_7255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7256 = {1{`RANDOM}};
  _T_3823_re = _RAND_7256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7257 = {1{`RANDOM}};
  _T_3823_im = _RAND_7257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7258 = {1{`RANDOM}};
  _T_3824_re = _RAND_7258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7259 = {1{`RANDOM}};
  _T_3824_im = _RAND_7259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7260 = {1{`RANDOM}};
  _T_3825_re = _RAND_7260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7261 = {1{`RANDOM}};
  _T_3825_im = _RAND_7261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7262 = {1{`RANDOM}};
  _T_3826_re = _RAND_7262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7263 = {1{`RANDOM}};
  _T_3826_im = _RAND_7263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7264 = {1{`RANDOM}};
  _T_3827_re = _RAND_7264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7265 = {1{`RANDOM}};
  _T_3827_im = _RAND_7265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7266 = {1{`RANDOM}};
  _T_3828_re = _RAND_7266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7267 = {1{`RANDOM}};
  _T_3828_im = _RAND_7267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7268 = {1{`RANDOM}};
  _T_3829_re = _RAND_7268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7269 = {1{`RANDOM}};
  _T_3829_im = _RAND_7269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7270 = {1{`RANDOM}};
  _T_3830_re = _RAND_7270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7271 = {1{`RANDOM}};
  _T_3830_im = _RAND_7271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7272 = {1{`RANDOM}};
  _T_3831_re = _RAND_7272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7273 = {1{`RANDOM}};
  _T_3831_im = _RAND_7273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7274 = {1{`RANDOM}};
  _T_3832_re = _RAND_7274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7275 = {1{`RANDOM}};
  _T_3832_im = _RAND_7275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7276 = {1{`RANDOM}};
  _T_3833_re = _RAND_7276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7277 = {1{`RANDOM}};
  _T_3833_im = _RAND_7277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7278 = {1{`RANDOM}};
  _T_3834_re = _RAND_7278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7279 = {1{`RANDOM}};
  _T_3834_im = _RAND_7279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7280 = {1{`RANDOM}};
  _T_3835_re = _RAND_7280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7281 = {1{`RANDOM}};
  _T_3835_im = _RAND_7281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7282 = {1{`RANDOM}};
  _T_3836_re = _RAND_7282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7283 = {1{`RANDOM}};
  _T_3836_im = _RAND_7283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7284 = {1{`RANDOM}};
  _T_3837_re = _RAND_7284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7285 = {1{`RANDOM}};
  _T_3837_im = _RAND_7285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7286 = {1{`RANDOM}};
  _T_3838_re = _RAND_7286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7287 = {1{`RANDOM}};
  _T_3838_im = _RAND_7287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7288 = {1{`RANDOM}};
  _T_3839_re = _RAND_7288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7289 = {1{`RANDOM}};
  _T_3839_im = _RAND_7289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7290 = {1{`RANDOM}};
  _T_3840_re = _RAND_7290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7291 = {1{`RANDOM}};
  _T_3840_im = _RAND_7291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7292 = {1{`RANDOM}};
  _T_3841_re = _RAND_7292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7293 = {1{`RANDOM}};
  _T_3841_im = _RAND_7293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7294 = {1{`RANDOM}};
  _T_3842_re = _RAND_7294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7295 = {1{`RANDOM}};
  _T_3842_im = _RAND_7295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7296 = {1{`RANDOM}};
  _T_3843_re = _RAND_7296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7297 = {1{`RANDOM}};
  _T_3843_im = _RAND_7297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7298 = {1{`RANDOM}};
  _T_3844_re = _RAND_7298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7299 = {1{`RANDOM}};
  _T_3844_im = _RAND_7299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7300 = {1{`RANDOM}};
  _T_3845_re = _RAND_7300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7301 = {1{`RANDOM}};
  _T_3845_im = _RAND_7301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7302 = {1{`RANDOM}};
  _T_3846_re = _RAND_7302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7303 = {1{`RANDOM}};
  _T_3846_im = _RAND_7303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7304 = {1{`RANDOM}};
  _T_3847_re = _RAND_7304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7305 = {1{`RANDOM}};
  _T_3847_im = _RAND_7305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7306 = {1{`RANDOM}};
  _T_3848_re = _RAND_7306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7307 = {1{`RANDOM}};
  _T_3848_im = _RAND_7307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7308 = {1{`RANDOM}};
  _T_3849_re = _RAND_7308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7309 = {1{`RANDOM}};
  _T_3849_im = _RAND_7309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7310 = {1{`RANDOM}};
  _T_3850_re = _RAND_7310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7311 = {1{`RANDOM}};
  _T_3850_im = _RAND_7311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7312 = {1{`RANDOM}};
  _T_3851_re = _RAND_7312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7313 = {1{`RANDOM}};
  _T_3851_im = _RAND_7313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7314 = {1{`RANDOM}};
  _T_3852_re = _RAND_7314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7315 = {1{`RANDOM}};
  _T_3852_im = _RAND_7315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7316 = {1{`RANDOM}};
  _T_3853_re = _RAND_7316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7317 = {1{`RANDOM}};
  _T_3853_im = _RAND_7317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7318 = {1{`RANDOM}};
  _T_3854_re = _RAND_7318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7319 = {1{`RANDOM}};
  _T_3854_im = _RAND_7319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7320 = {1{`RANDOM}};
  _T_3855_re = _RAND_7320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7321 = {1{`RANDOM}};
  _T_3855_im = _RAND_7321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7322 = {1{`RANDOM}};
  _T_3856_re = _RAND_7322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7323 = {1{`RANDOM}};
  _T_3856_im = _RAND_7323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7324 = {1{`RANDOM}};
  _T_3857_re = _RAND_7324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7325 = {1{`RANDOM}};
  _T_3857_im = _RAND_7325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7326 = {1{`RANDOM}};
  _T_3858_re = _RAND_7326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7327 = {1{`RANDOM}};
  _T_3858_im = _RAND_7327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7328 = {1{`RANDOM}};
  _T_3859_re = _RAND_7328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7329 = {1{`RANDOM}};
  _T_3859_im = _RAND_7329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7330 = {1{`RANDOM}};
  _T_3860_re = _RAND_7330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7331 = {1{`RANDOM}};
  _T_3860_im = _RAND_7331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7332 = {1{`RANDOM}};
  _T_3861_re = _RAND_7332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7333 = {1{`RANDOM}};
  _T_3861_im = _RAND_7333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7334 = {1{`RANDOM}};
  _T_3862_re = _RAND_7334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7335 = {1{`RANDOM}};
  _T_3862_im = _RAND_7335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7336 = {1{`RANDOM}};
  _T_3863_re = _RAND_7336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7337 = {1{`RANDOM}};
  _T_3863_im = _RAND_7337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7338 = {1{`RANDOM}};
  _T_3864_re = _RAND_7338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7339 = {1{`RANDOM}};
  _T_3864_im = _RAND_7339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7340 = {1{`RANDOM}};
  _T_3865_re = _RAND_7340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7341 = {1{`RANDOM}};
  _T_3865_im = _RAND_7341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7342 = {1{`RANDOM}};
  _T_3866_re = _RAND_7342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7343 = {1{`RANDOM}};
  _T_3866_im = _RAND_7343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7344 = {1{`RANDOM}};
  _T_3867_re = _RAND_7344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7345 = {1{`RANDOM}};
  _T_3867_im = _RAND_7345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7346 = {1{`RANDOM}};
  _T_3868_re = _RAND_7346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7347 = {1{`RANDOM}};
  _T_3868_im = _RAND_7347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7348 = {1{`RANDOM}};
  _T_3869_re = _RAND_7348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7349 = {1{`RANDOM}};
  _T_3869_im = _RAND_7349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7350 = {1{`RANDOM}};
  _T_3870_re = _RAND_7350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7351 = {1{`RANDOM}};
  _T_3870_im = _RAND_7351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7352 = {1{`RANDOM}};
  _T_3871_re = _RAND_7352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7353 = {1{`RANDOM}};
  _T_3871_im = _RAND_7353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7354 = {1{`RANDOM}};
  _T_3872_re = _RAND_7354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7355 = {1{`RANDOM}};
  _T_3872_im = _RAND_7355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7356 = {1{`RANDOM}};
  _T_3873_re = _RAND_7356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7357 = {1{`RANDOM}};
  _T_3873_im = _RAND_7357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7358 = {1{`RANDOM}};
  _T_3874_re = _RAND_7358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7359 = {1{`RANDOM}};
  _T_3874_im = _RAND_7359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7360 = {1{`RANDOM}};
  _T_3875_re = _RAND_7360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7361 = {1{`RANDOM}};
  _T_3875_im = _RAND_7361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7362 = {1{`RANDOM}};
  _T_3876_re = _RAND_7362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7363 = {1{`RANDOM}};
  _T_3876_im = _RAND_7363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7364 = {1{`RANDOM}};
  _T_3877_re = _RAND_7364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7365 = {1{`RANDOM}};
  _T_3877_im = _RAND_7365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7366 = {1{`RANDOM}};
  _T_3878_re = _RAND_7366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7367 = {1{`RANDOM}};
  _T_3878_im = _RAND_7367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7368 = {1{`RANDOM}};
  _T_3879_re = _RAND_7368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7369 = {1{`RANDOM}};
  _T_3879_im = _RAND_7369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7370 = {1{`RANDOM}};
  _T_3880_re = _RAND_7370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7371 = {1{`RANDOM}};
  _T_3880_im = _RAND_7371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7372 = {1{`RANDOM}};
  _T_3881_re = _RAND_7372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7373 = {1{`RANDOM}};
  _T_3881_im = _RAND_7373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7374 = {1{`RANDOM}};
  _T_3882_re = _RAND_7374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7375 = {1{`RANDOM}};
  _T_3882_im = _RAND_7375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7376 = {1{`RANDOM}};
  _T_3883_re = _RAND_7376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7377 = {1{`RANDOM}};
  _T_3883_im = _RAND_7377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7378 = {1{`RANDOM}};
  _T_3884_re = _RAND_7378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7379 = {1{`RANDOM}};
  _T_3884_im = _RAND_7379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7380 = {1{`RANDOM}};
  _T_3885_re = _RAND_7380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7381 = {1{`RANDOM}};
  _T_3885_im = _RAND_7381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7382 = {1{`RANDOM}};
  _T_3886_re = _RAND_7382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7383 = {1{`RANDOM}};
  _T_3886_im = _RAND_7383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7384 = {1{`RANDOM}};
  _T_3887_re = _RAND_7384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7385 = {1{`RANDOM}};
  _T_3887_im = _RAND_7385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7386 = {1{`RANDOM}};
  _T_3888_re = _RAND_7386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7387 = {1{`RANDOM}};
  _T_3888_im = _RAND_7387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7388 = {1{`RANDOM}};
  _T_3889_re = _RAND_7388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7389 = {1{`RANDOM}};
  _T_3889_im = _RAND_7389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7390 = {1{`RANDOM}};
  _T_3890_re = _RAND_7390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7391 = {1{`RANDOM}};
  _T_3890_im = _RAND_7391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7392 = {1{`RANDOM}};
  _T_3891_re = _RAND_7392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7393 = {1{`RANDOM}};
  _T_3891_im = _RAND_7393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7394 = {1{`RANDOM}};
  _T_3892_re = _RAND_7394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7395 = {1{`RANDOM}};
  _T_3892_im = _RAND_7395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7396 = {1{`RANDOM}};
  _T_3893_re = _RAND_7396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7397 = {1{`RANDOM}};
  _T_3893_im = _RAND_7397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7398 = {1{`RANDOM}};
  _T_3894_re = _RAND_7398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7399 = {1{`RANDOM}};
  _T_3894_im = _RAND_7399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7400 = {1{`RANDOM}};
  _T_3895_re = _RAND_7400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7401 = {1{`RANDOM}};
  _T_3895_im = _RAND_7401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7402 = {1{`RANDOM}};
  _T_3896_re = _RAND_7402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7403 = {1{`RANDOM}};
  _T_3896_im = _RAND_7403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7404 = {1{`RANDOM}};
  _T_3897_re = _RAND_7404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7405 = {1{`RANDOM}};
  _T_3897_im = _RAND_7405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7406 = {1{`RANDOM}};
  _T_3898_re = _RAND_7406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7407 = {1{`RANDOM}};
  _T_3898_im = _RAND_7407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7408 = {1{`RANDOM}};
  _T_3899_re = _RAND_7408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7409 = {1{`RANDOM}};
  _T_3899_im = _RAND_7409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7410 = {1{`RANDOM}};
  _T_3900_re = _RAND_7410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7411 = {1{`RANDOM}};
  _T_3900_im = _RAND_7411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7412 = {1{`RANDOM}};
  _T_3901_re = _RAND_7412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7413 = {1{`RANDOM}};
  _T_3901_im = _RAND_7413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7414 = {1{`RANDOM}};
  _T_3902_re = _RAND_7414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7415 = {1{`RANDOM}};
  _T_3902_im = _RAND_7415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7416 = {1{`RANDOM}};
  _T_3903_re = _RAND_7416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7417 = {1{`RANDOM}};
  _T_3903_im = _RAND_7417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7418 = {1{`RANDOM}};
  _T_3904_re = _RAND_7418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7419 = {1{`RANDOM}};
  _T_3904_im = _RAND_7419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7420 = {1{`RANDOM}};
  _T_3905_re = _RAND_7420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7421 = {1{`RANDOM}};
  _T_3905_im = _RAND_7421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7422 = {1{`RANDOM}};
  _T_3906_re = _RAND_7422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7423 = {1{`RANDOM}};
  _T_3906_im = _RAND_7423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7424 = {1{`RANDOM}};
  _T_3907_re = _RAND_7424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7425 = {1{`RANDOM}};
  _T_3907_im = _RAND_7425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7426 = {1{`RANDOM}};
  _T_3908_re = _RAND_7426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7427 = {1{`RANDOM}};
  _T_3908_im = _RAND_7427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7428 = {1{`RANDOM}};
  _T_3909_re = _RAND_7428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7429 = {1{`RANDOM}};
  _T_3909_im = _RAND_7429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7430 = {1{`RANDOM}};
  _T_3910_re = _RAND_7430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7431 = {1{`RANDOM}};
  _T_3910_im = _RAND_7431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7432 = {1{`RANDOM}};
  _T_3911_re = _RAND_7432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7433 = {1{`RANDOM}};
  _T_3911_im = _RAND_7433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7434 = {1{`RANDOM}};
  _T_3912_re = _RAND_7434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7435 = {1{`RANDOM}};
  _T_3912_im = _RAND_7435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7436 = {1{`RANDOM}};
  _T_3913_re = _RAND_7436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7437 = {1{`RANDOM}};
  _T_3913_im = _RAND_7437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7438 = {1{`RANDOM}};
  _T_3914_re = _RAND_7438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7439 = {1{`RANDOM}};
  _T_3914_im = _RAND_7439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7440 = {1{`RANDOM}};
  _T_3915_re = _RAND_7440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7441 = {1{`RANDOM}};
  _T_3915_im = _RAND_7441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7442 = {1{`RANDOM}};
  _T_3916_re = _RAND_7442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7443 = {1{`RANDOM}};
  _T_3916_im = _RAND_7443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7444 = {1{`RANDOM}};
  _T_3917_re = _RAND_7444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7445 = {1{`RANDOM}};
  _T_3917_im = _RAND_7445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7446 = {1{`RANDOM}};
  _T_3918_re = _RAND_7446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7447 = {1{`RANDOM}};
  _T_3918_im = _RAND_7447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7448 = {1{`RANDOM}};
  _T_3919_re = _RAND_7448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7449 = {1{`RANDOM}};
  _T_3919_im = _RAND_7449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7450 = {1{`RANDOM}};
  _T_3920_re = _RAND_7450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7451 = {1{`RANDOM}};
  _T_3920_im = _RAND_7451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7452 = {1{`RANDOM}};
  _T_3921_re = _RAND_7452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7453 = {1{`RANDOM}};
  _T_3921_im = _RAND_7453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7454 = {1{`RANDOM}};
  _T_3922_re = _RAND_7454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7455 = {1{`RANDOM}};
  _T_3922_im = _RAND_7455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7456 = {1{`RANDOM}};
  _T_3923_re = _RAND_7456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7457 = {1{`RANDOM}};
  _T_3923_im = _RAND_7457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7458 = {1{`RANDOM}};
  _T_3924_re = _RAND_7458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7459 = {1{`RANDOM}};
  _T_3924_im = _RAND_7459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7460 = {1{`RANDOM}};
  _T_3925_re = _RAND_7460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7461 = {1{`RANDOM}};
  _T_3925_im = _RAND_7461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7462 = {1{`RANDOM}};
  _T_3926_re = _RAND_7462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7463 = {1{`RANDOM}};
  _T_3926_im = _RAND_7463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7464 = {1{`RANDOM}};
  _T_3927_re = _RAND_7464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7465 = {1{`RANDOM}};
  _T_3927_im = _RAND_7465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7466 = {1{`RANDOM}};
  _T_3928_re = _RAND_7466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7467 = {1{`RANDOM}};
  _T_3928_im = _RAND_7467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7468 = {1{`RANDOM}};
  _T_3929_re = _RAND_7468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7469 = {1{`RANDOM}};
  _T_3929_im = _RAND_7469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7470 = {1{`RANDOM}};
  _T_3930_re = _RAND_7470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7471 = {1{`RANDOM}};
  _T_3930_im = _RAND_7471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7472 = {1{`RANDOM}};
  _T_3931_re = _RAND_7472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7473 = {1{`RANDOM}};
  _T_3931_im = _RAND_7473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7474 = {1{`RANDOM}};
  _T_3932_re = _RAND_7474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7475 = {1{`RANDOM}};
  _T_3932_im = _RAND_7475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7476 = {1{`RANDOM}};
  _T_3933_re = _RAND_7476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7477 = {1{`RANDOM}};
  _T_3933_im = _RAND_7477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7478 = {1{`RANDOM}};
  _T_3934_re = _RAND_7478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7479 = {1{`RANDOM}};
  _T_3934_im = _RAND_7479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7480 = {1{`RANDOM}};
  _T_3935_re = _RAND_7480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7481 = {1{`RANDOM}};
  _T_3935_im = _RAND_7481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7482 = {1{`RANDOM}};
  _T_3936_re = _RAND_7482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7483 = {1{`RANDOM}};
  _T_3936_im = _RAND_7483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7484 = {1{`RANDOM}};
  _T_3937_re = _RAND_7484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7485 = {1{`RANDOM}};
  _T_3937_im = _RAND_7485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7486 = {1{`RANDOM}};
  _T_3938_re = _RAND_7486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7487 = {1{`RANDOM}};
  _T_3938_im = _RAND_7487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7488 = {1{`RANDOM}};
  _T_3939_re = _RAND_7488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7489 = {1{`RANDOM}};
  _T_3939_im = _RAND_7489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7490 = {1{`RANDOM}};
  _T_3940_re = _RAND_7490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7491 = {1{`RANDOM}};
  _T_3940_im = _RAND_7491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7492 = {1{`RANDOM}};
  _T_3941_re = _RAND_7492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7493 = {1{`RANDOM}};
  _T_3941_im = _RAND_7493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7494 = {1{`RANDOM}};
  _T_3942_re = _RAND_7494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7495 = {1{`RANDOM}};
  _T_3942_im = _RAND_7495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7496 = {1{`RANDOM}};
  _T_3943_re = _RAND_7496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7497 = {1{`RANDOM}};
  _T_3943_im = _RAND_7497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7498 = {1{`RANDOM}};
  _T_3944_re = _RAND_7498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7499 = {1{`RANDOM}};
  _T_3944_im = _RAND_7499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7500 = {1{`RANDOM}};
  _T_3945_re = _RAND_7500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7501 = {1{`RANDOM}};
  _T_3945_im = _RAND_7501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7502 = {1{`RANDOM}};
  _T_3946_re = _RAND_7502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7503 = {1{`RANDOM}};
  _T_3946_im = _RAND_7503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7504 = {1{`RANDOM}};
  _T_3947_re = _RAND_7504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7505 = {1{`RANDOM}};
  _T_3947_im = _RAND_7505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7506 = {1{`RANDOM}};
  _T_3948_re = _RAND_7506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7507 = {1{`RANDOM}};
  _T_3948_im = _RAND_7507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7508 = {1{`RANDOM}};
  _T_3949_re = _RAND_7508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7509 = {1{`RANDOM}};
  _T_3949_im = _RAND_7509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7510 = {1{`RANDOM}};
  _T_3950_re = _RAND_7510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7511 = {1{`RANDOM}};
  _T_3950_im = _RAND_7511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7512 = {1{`RANDOM}};
  _T_3951_re = _RAND_7512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7513 = {1{`RANDOM}};
  _T_3951_im = _RAND_7513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7514 = {1{`RANDOM}};
  _T_3952_re = _RAND_7514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7515 = {1{`RANDOM}};
  _T_3952_im = _RAND_7515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7516 = {1{`RANDOM}};
  _T_3953_re = _RAND_7516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7517 = {1{`RANDOM}};
  _T_3953_im = _RAND_7517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7518 = {1{`RANDOM}};
  _T_3954_re = _RAND_7518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7519 = {1{`RANDOM}};
  _T_3954_im = _RAND_7519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7520 = {1{`RANDOM}};
  _T_3955_re = _RAND_7520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7521 = {1{`RANDOM}};
  _T_3955_im = _RAND_7521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7522 = {1{`RANDOM}};
  _T_3956_re = _RAND_7522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7523 = {1{`RANDOM}};
  _T_3956_im = _RAND_7523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7524 = {1{`RANDOM}};
  _T_3957_re = _RAND_7524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7525 = {1{`RANDOM}};
  _T_3957_im = _RAND_7525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7526 = {1{`RANDOM}};
  _T_3958_re = _RAND_7526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7527 = {1{`RANDOM}};
  _T_3958_im = _RAND_7527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7528 = {1{`RANDOM}};
  _T_3959_re = _RAND_7528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7529 = {1{`RANDOM}};
  _T_3959_im = _RAND_7529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7530 = {1{`RANDOM}};
  _T_3960_re = _RAND_7530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7531 = {1{`RANDOM}};
  _T_3960_im = _RAND_7531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7532 = {1{`RANDOM}};
  _T_3961_re = _RAND_7532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7533 = {1{`RANDOM}};
  _T_3961_im = _RAND_7533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7534 = {1{`RANDOM}};
  _T_3962_re = _RAND_7534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7535 = {1{`RANDOM}};
  _T_3962_im = _RAND_7535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7536 = {1{`RANDOM}};
  _T_3963_re = _RAND_7536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7537 = {1{`RANDOM}};
  _T_3963_im = _RAND_7537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7538 = {1{`RANDOM}};
  _T_3964_re = _RAND_7538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7539 = {1{`RANDOM}};
  _T_3964_im = _RAND_7539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7540 = {1{`RANDOM}};
  _T_3965_re = _RAND_7540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7541 = {1{`RANDOM}};
  _T_3965_im = _RAND_7541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7542 = {1{`RANDOM}};
  _T_3966_re = _RAND_7542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7543 = {1{`RANDOM}};
  _T_3966_im = _RAND_7543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7544 = {1{`RANDOM}};
  _T_3967_re = _RAND_7544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7545 = {1{`RANDOM}};
  _T_3967_im = _RAND_7545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7546 = {1{`RANDOM}};
  _T_3968_re = _RAND_7546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7547 = {1{`RANDOM}};
  _T_3968_im = _RAND_7547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7548 = {1{`RANDOM}};
  _T_3969_re = _RAND_7548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7549 = {1{`RANDOM}};
  _T_3969_im = _RAND_7549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7550 = {1{`RANDOM}};
  _T_3970_re = _RAND_7550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7551 = {1{`RANDOM}};
  _T_3970_im = _RAND_7551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7552 = {1{`RANDOM}};
  _T_3971_re = _RAND_7552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7553 = {1{`RANDOM}};
  _T_3971_im = _RAND_7553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7554 = {1{`RANDOM}};
  _T_3972_re = _RAND_7554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7555 = {1{`RANDOM}};
  _T_3972_im = _RAND_7555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7556 = {1{`RANDOM}};
  _T_3973_re = _RAND_7556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7557 = {1{`RANDOM}};
  _T_3973_im = _RAND_7557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7558 = {1{`RANDOM}};
  _T_3974_re = _RAND_7558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7559 = {1{`RANDOM}};
  _T_3974_im = _RAND_7559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7560 = {1{`RANDOM}};
  _T_3975_re = _RAND_7560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7561 = {1{`RANDOM}};
  _T_3975_im = _RAND_7561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7562 = {1{`RANDOM}};
  _T_3976_re = _RAND_7562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7563 = {1{`RANDOM}};
  _T_3976_im = _RAND_7563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7564 = {1{`RANDOM}};
  _T_3977_re = _RAND_7564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7565 = {1{`RANDOM}};
  _T_3977_im = _RAND_7565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7566 = {1{`RANDOM}};
  _T_3978_re = _RAND_7566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7567 = {1{`RANDOM}};
  _T_3978_im = _RAND_7567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7568 = {1{`RANDOM}};
  _T_3979_re = _RAND_7568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7569 = {1{`RANDOM}};
  _T_3979_im = _RAND_7569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7570 = {1{`RANDOM}};
  _T_3980_re = _RAND_7570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7571 = {1{`RANDOM}};
  _T_3980_im = _RAND_7571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7572 = {1{`RANDOM}};
  _T_3981_re = _RAND_7572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7573 = {1{`RANDOM}};
  _T_3981_im = _RAND_7573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7574 = {1{`RANDOM}};
  _T_3982_re = _RAND_7574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7575 = {1{`RANDOM}};
  _T_3982_im = _RAND_7575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7576 = {1{`RANDOM}};
  _T_3983_re = _RAND_7576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7577 = {1{`RANDOM}};
  _T_3983_im = _RAND_7577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7578 = {1{`RANDOM}};
  _T_3984_re = _RAND_7578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7579 = {1{`RANDOM}};
  _T_3984_im = _RAND_7579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7580 = {1{`RANDOM}};
  _T_3985_re = _RAND_7580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7581 = {1{`RANDOM}};
  _T_3985_im = _RAND_7581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7582 = {1{`RANDOM}};
  _T_3986_re = _RAND_7582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7583 = {1{`RANDOM}};
  _T_3986_im = _RAND_7583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7584 = {1{`RANDOM}};
  _T_3987_re = _RAND_7584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7585 = {1{`RANDOM}};
  _T_3987_im = _RAND_7585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7586 = {1{`RANDOM}};
  _T_3988_re = _RAND_7586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7587 = {1{`RANDOM}};
  _T_3988_im = _RAND_7587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7588 = {1{`RANDOM}};
  _T_3989_re = _RAND_7588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7589 = {1{`RANDOM}};
  _T_3989_im = _RAND_7589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7590 = {1{`RANDOM}};
  _T_3990_re = _RAND_7590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7591 = {1{`RANDOM}};
  _T_3990_im = _RAND_7591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7592 = {1{`RANDOM}};
  _T_3991_re = _RAND_7592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7593 = {1{`RANDOM}};
  _T_3991_im = _RAND_7593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7594 = {1{`RANDOM}};
  _T_3992_re = _RAND_7594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7595 = {1{`RANDOM}};
  _T_3992_im = _RAND_7595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7596 = {1{`RANDOM}};
  _T_3993_re = _RAND_7596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7597 = {1{`RANDOM}};
  _T_3993_im = _RAND_7597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7598 = {1{`RANDOM}};
  _T_3994_re = _RAND_7598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7599 = {1{`RANDOM}};
  _T_3994_im = _RAND_7599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7600 = {1{`RANDOM}};
  _T_3995_re = _RAND_7600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7601 = {1{`RANDOM}};
  _T_3995_im = _RAND_7601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7602 = {1{`RANDOM}};
  _T_3996_re = _RAND_7602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7603 = {1{`RANDOM}};
  _T_3996_im = _RAND_7603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7604 = {1{`RANDOM}};
  _T_3997_re = _RAND_7604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7605 = {1{`RANDOM}};
  _T_3997_im = _RAND_7605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7606 = {1{`RANDOM}};
  _T_3998_re = _RAND_7606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7607 = {1{`RANDOM}};
  _T_3998_im = _RAND_7607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7608 = {1{`RANDOM}};
  _T_3999_re = _RAND_7608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7609 = {1{`RANDOM}};
  _T_3999_im = _RAND_7609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7610 = {1{`RANDOM}};
  _T_4000_re = _RAND_7610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7611 = {1{`RANDOM}};
  _T_4000_im = _RAND_7611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7612 = {1{`RANDOM}};
  _T_4001_re = _RAND_7612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7613 = {1{`RANDOM}};
  _T_4001_im = _RAND_7613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7614 = {1{`RANDOM}};
  _T_4002_re = _RAND_7614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7615 = {1{`RANDOM}};
  _T_4002_im = _RAND_7615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7616 = {1{`RANDOM}};
  _T_4003_re = _RAND_7616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7617 = {1{`RANDOM}};
  _T_4003_im = _RAND_7617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7618 = {1{`RANDOM}};
  _T_4004_re = _RAND_7618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7619 = {1{`RANDOM}};
  _T_4004_im = _RAND_7619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7620 = {1{`RANDOM}};
  _T_4005_re = _RAND_7620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7621 = {1{`RANDOM}};
  _T_4005_im = _RAND_7621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7622 = {1{`RANDOM}};
  _T_4006_re = _RAND_7622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7623 = {1{`RANDOM}};
  _T_4006_im = _RAND_7623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7624 = {1{`RANDOM}};
  _T_4007_re = _RAND_7624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7625 = {1{`RANDOM}};
  _T_4007_im = _RAND_7625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7626 = {1{`RANDOM}};
  _T_4008_re = _RAND_7626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7627 = {1{`RANDOM}};
  _T_4008_im = _RAND_7627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7628 = {1{`RANDOM}};
  _T_4009_re = _RAND_7628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7629 = {1{`RANDOM}};
  _T_4009_im = _RAND_7629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7630 = {1{`RANDOM}};
  _T_4010_re = _RAND_7630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7631 = {1{`RANDOM}};
  _T_4010_im = _RAND_7631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7632 = {1{`RANDOM}};
  _T_4011_re = _RAND_7632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7633 = {1{`RANDOM}};
  _T_4011_im = _RAND_7633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7634 = {1{`RANDOM}};
  _T_4012_re = _RAND_7634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7635 = {1{`RANDOM}};
  _T_4012_im = _RAND_7635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7636 = {1{`RANDOM}};
  _T_4013_re = _RAND_7636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7637 = {1{`RANDOM}};
  _T_4013_im = _RAND_7637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7638 = {1{`RANDOM}};
  _T_4014_re = _RAND_7638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7639 = {1{`RANDOM}};
  _T_4014_im = _RAND_7639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7640 = {1{`RANDOM}};
  _T_4015_re = _RAND_7640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7641 = {1{`RANDOM}};
  _T_4015_im = _RAND_7641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7642 = {1{`RANDOM}};
  _T_4016_re = _RAND_7642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7643 = {1{`RANDOM}};
  _T_4016_im = _RAND_7643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7644 = {1{`RANDOM}};
  _T_4017_re = _RAND_7644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7645 = {1{`RANDOM}};
  _T_4017_im = _RAND_7645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7646 = {1{`RANDOM}};
  _T_4018_re = _RAND_7646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7647 = {1{`RANDOM}};
  _T_4018_im = _RAND_7647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7648 = {1{`RANDOM}};
  _T_4019_re = _RAND_7648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7649 = {1{`RANDOM}};
  _T_4019_im = _RAND_7649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7650 = {1{`RANDOM}};
  _T_4020_re = _RAND_7650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7651 = {1{`RANDOM}};
  _T_4020_im = _RAND_7651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7652 = {1{`RANDOM}};
  _T_4021_re = _RAND_7652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7653 = {1{`RANDOM}};
  _T_4021_im = _RAND_7653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7654 = {1{`RANDOM}};
  _T_4022_re = _RAND_7654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7655 = {1{`RANDOM}};
  _T_4022_im = _RAND_7655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7656 = {1{`RANDOM}};
  _T_4023_re = _RAND_7656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7657 = {1{`RANDOM}};
  _T_4023_im = _RAND_7657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7658 = {1{`RANDOM}};
  _T_4024_re = _RAND_7658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7659 = {1{`RANDOM}};
  _T_4024_im = _RAND_7659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7660 = {1{`RANDOM}};
  _T_4025_re = _RAND_7660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7661 = {1{`RANDOM}};
  _T_4025_im = _RAND_7661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7662 = {1{`RANDOM}};
  _T_4026_re = _RAND_7662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7663 = {1{`RANDOM}};
  _T_4026_im = _RAND_7663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7664 = {1{`RANDOM}};
  _T_4027_re = _RAND_7664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7665 = {1{`RANDOM}};
  _T_4027_im = _RAND_7665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7666 = {1{`RANDOM}};
  _T_4028_re = _RAND_7666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7667 = {1{`RANDOM}};
  _T_4028_im = _RAND_7667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7668 = {1{`RANDOM}};
  _T_4029_re = _RAND_7668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7669 = {1{`RANDOM}};
  _T_4029_im = _RAND_7669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7670 = {1{`RANDOM}};
  _T_4030_re = _RAND_7670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7671 = {1{`RANDOM}};
  _T_4030_im = _RAND_7671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7672 = {1{`RANDOM}};
  _T_4031_re = _RAND_7672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7673 = {1{`RANDOM}};
  _T_4031_im = _RAND_7673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7674 = {1{`RANDOM}};
  _T_4032_re = _RAND_7674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7675 = {1{`RANDOM}};
  _T_4032_im = _RAND_7675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7676 = {1{`RANDOM}};
  _T_4033_re = _RAND_7676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7677 = {1{`RANDOM}};
  _T_4033_im = _RAND_7677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7678 = {1{`RANDOM}};
  _T_4034_re = _RAND_7678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7679 = {1{`RANDOM}};
  _T_4034_im = _RAND_7679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7680 = {1{`RANDOM}};
  _T_4035_re = _RAND_7680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7681 = {1{`RANDOM}};
  _T_4035_im = _RAND_7681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7682 = {1{`RANDOM}};
  _T_4036_re = _RAND_7682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7683 = {1{`RANDOM}};
  _T_4036_im = _RAND_7683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7684 = {1{`RANDOM}};
  _T_4037_re = _RAND_7684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7685 = {1{`RANDOM}};
  _T_4037_im = _RAND_7685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7686 = {1{`RANDOM}};
  _T_4038_re = _RAND_7686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7687 = {1{`RANDOM}};
  _T_4038_im = _RAND_7687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7688 = {1{`RANDOM}};
  _T_4039_re = _RAND_7688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7689 = {1{`RANDOM}};
  _T_4039_im = _RAND_7689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7690 = {1{`RANDOM}};
  _T_4040_re = _RAND_7690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7691 = {1{`RANDOM}};
  _T_4040_im = _RAND_7691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7692 = {1{`RANDOM}};
  _T_4041_re = _RAND_7692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7693 = {1{`RANDOM}};
  _T_4041_im = _RAND_7693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7694 = {1{`RANDOM}};
  _T_4042_re = _RAND_7694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7695 = {1{`RANDOM}};
  _T_4042_im = _RAND_7695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7696 = {1{`RANDOM}};
  _T_4043_re = _RAND_7696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7697 = {1{`RANDOM}};
  _T_4043_im = _RAND_7697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7698 = {1{`RANDOM}};
  _T_4044_re = _RAND_7698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7699 = {1{`RANDOM}};
  _T_4044_im = _RAND_7699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7700 = {1{`RANDOM}};
  _T_4045_re = _RAND_7700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7701 = {1{`RANDOM}};
  _T_4045_im = _RAND_7701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7702 = {1{`RANDOM}};
  _T_4046_re = _RAND_7702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7703 = {1{`RANDOM}};
  _T_4046_im = _RAND_7703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7704 = {1{`RANDOM}};
  _T_4047_re = _RAND_7704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7705 = {1{`RANDOM}};
  _T_4047_im = _RAND_7705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7706 = {1{`RANDOM}};
  _T_4048_re = _RAND_7706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7707 = {1{`RANDOM}};
  _T_4048_im = _RAND_7707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7708 = {1{`RANDOM}};
  _T_4049_re = _RAND_7708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7709 = {1{`RANDOM}};
  _T_4049_im = _RAND_7709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7710 = {1{`RANDOM}};
  _T_4050_re = _RAND_7710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7711 = {1{`RANDOM}};
  _T_4050_im = _RAND_7711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7712 = {1{`RANDOM}};
  _T_4051_re = _RAND_7712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7713 = {1{`RANDOM}};
  _T_4051_im = _RAND_7713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7714 = {1{`RANDOM}};
  _T_4052_re = _RAND_7714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7715 = {1{`RANDOM}};
  _T_4052_im = _RAND_7715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7716 = {1{`RANDOM}};
  _T_4053_re = _RAND_7716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7717 = {1{`RANDOM}};
  _T_4053_im = _RAND_7717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7718 = {1{`RANDOM}};
  _T_4054_re = _RAND_7718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7719 = {1{`RANDOM}};
  _T_4054_im = _RAND_7719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7720 = {1{`RANDOM}};
  _T_4055_re = _RAND_7720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7721 = {1{`RANDOM}};
  _T_4055_im = _RAND_7721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7722 = {1{`RANDOM}};
  _T_4056_re = _RAND_7722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7723 = {1{`RANDOM}};
  _T_4056_im = _RAND_7723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7724 = {1{`RANDOM}};
  _T_4057_re = _RAND_7724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7725 = {1{`RANDOM}};
  _T_4057_im = _RAND_7725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7726 = {1{`RANDOM}};
  _T_4058_re = _RAND_7726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7727 = {1{`RANDOM}};
  _T_4058_im = _RAND_7727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7728 = {1{`RANDOM}};
  _T_4059_re = _RAND_7728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7729 = {1{`RANDOM}};
  _T_4059_im = _RAND_7729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7730 = {1{`RANDOM}};
  _T_4060_re = _RAND_7730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7731 = {1{`RANDOM}};
  _T_4060_im = _RAND_7731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7732 = {1{`RANDOM}};
  _T_4061_re = _RAND_7732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7733 = {1{`RANDOM}};
  _T_4061_im = _RAND_7733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7734 = {1{`RANDOM}};
  _T_4062_re = _RAND_7734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7735 = {1{`RANDOM}};
  _T_4062_im = _RAND_7735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7736 = {1{`RANDOM}};
  _T_4063_re = _RAND_7736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7737 = {1{`RANDOM}};
  _T_4063_im = _RAND_7737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7738 = {1{`RANDOM}};
  _T_4064_re = _RAND_7738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7739 = {1{`RANDOM}};
  _T_4064_im = _RAND_7739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7740 = {1{`RANDOM}};
  _T_4065_re = _RAND_7740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7741 = {1{`RANDOM}};
  _T_4065_im = _RAND_7741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7742 = {1{`RANDOM}};
  _T_4066_re = _RAND_7742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7743 = {1{`RANDOM}};
  _T_4066_im = _RAND_7743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7744 = {1{`RANDOM}};
  _T_4067_re = _RAND_7744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7745 = {1{`RANDOM}};
  _T_4067_im = _RAND_7745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7746 = {1{`RANDOM}};
  _T_4068_re = _RAND_7746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7747 = {1{`RANDOM}};
  _T_4068_im = _RAND_7747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7748 = {1{`RANDOM}};
  _T_4069_re = _RAND_7748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7749 = {1{`RANDOM}};
  _T_4069_im = _RAND_7749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7750 = {1{`RANDOM}};
  _T_4070_re = _RAND_7750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7751 = {1{`RANDOM}};
  _T_4070_im = _RAND_7751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7752 = {1{`RANDOM}};
  _T_4071_re = _RAND_7752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7753 = {1{`RANDOM}};
  _T_4071_im = _RAND_7753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7754 = {1{`RANDOM}};
  _T_4072_re = _RAND_7754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7755 = {1{`RANDOM}};
  _T_4072_im = _RAND_7755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7756 = {1{`RANDOM}};
  _T_4073_re = _RAND_7756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7757 = {1{`RANDOM}};
  _T_4073_im = _RAND_7757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7758 = {1{`RANDOM}};
  _T_4074_re = _RAND_7758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7759 = {1{`RANDOM}};
  _T_4074_im = _RAND_7759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7760 = {1{`RANDOM}};
  _T_4075_re = _RAND_7760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7761 = {1{`RANDOM}};
  _T_4075_im = _RAND_7761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7762 = {1{`RANDOM}};
  _T_4076_re = _RAND_7762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7763 = {1{`RANDOM}};
  _T_4076_im = _RAND_7763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7764 = {1{`RANDOM}};
  _T_4077_re = _RAND_7764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7765 = {1{`RANDOM}};
  _T_4077_im = _RAND_7765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7766 = {1{`RANDOM}};
  _T_4078_re = _RAND_7766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7767 = {1{`RANDOM}};
  _T_4078_im = _RAND_7767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7768 = {1{`RANDOM}};
  _T_4079_re = _RAND_7768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7769 = {1{`RANDOM}};
  _T_4079_im = _RAND_7769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7770 = {1{`RANDOM}};
  _T_4080_re = _RAND_7770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7771 = {1{`RANDOM}};
  _T_4080_im = _RAND_7771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7772 = {1{`RANDOM}};
  _T_4081_re = _RAND_7772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7773 = {1{`RANDOM}};
  _T_4081_im = _RAND_7773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7774 = {1{`RANDOM}};
  _T_4082_re = _RAND_7774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7775 = {1{`RANDOM}};
  _T_4082_im = _RAND_7775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7776 = {1{`RANDOM}};
  _T_4083_re = _RAND_7776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7777 = {1{`RANDOM}};
  _T_4083_im = _RAND_7777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7778 = {1{`RANDOM}};
  _T_4084_re = _RAND_7778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7779 = {1{`RANDOM}};
  _T_4084_im = _RAND_7779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7780 = {1{`RANDOM}};
  _T_4085_re = _RAND_7780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7781 = {1{`RANDOM}};
  _T_4085_im = _RAND_7781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7782 = {1{`RANDOM}};
  _T_4086_re = _RAND_7782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7783 = {1{`RANDOM}};
  _T_4086_im = _RAND_7783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7784 = {1{`RANDOM}};
  _T_4087_re = _RAND_7784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7785 = {1{`RANDOM}};
  _T_4087_im = _RAND_7785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7786 = {1{`RANDOM}};
  _T_4088_re = _RAND_7786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7787 = {1{`RANDOM}};
  _T_4088_im = _RAND_7787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7788 = {1{`RANDOM}};
  _T_4089_re = _RAND_7788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7789 = {1{`RANDOM}};
  _T_4089_im = _RAND_7789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7790 = {1{`RANDOM}};
  _T_4090_re = _RAND_7790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7791 = {1{`RANDOM}};
  _T_4090_im = _RAND_7791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7792 = {1{`RANDOM}};
  _T_4091_re = _RAND_7792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7793 = {1{`RANDOM}};
  _T_4091_im = _RAND_7793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7794 = {1{`RANDOM}};
  _T_4092_re = _RAND_7794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7795 = {1{`RANDOM}};
  _T_4092_im = _RAND_7795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7796 = {1{`RANDOM}};
  _T_4093_re = _RAND_7796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7797 = {1{`RANDOM}};
  _T_4093_im = _RAND_7797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7798 = {1{`RANDOM}};
  _T_4094_re = _RAND_7798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7799 = {1{`RANDOM}};
  _T_4094_im = _RAND_7799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7800 = {1{`RANDOM}};
  _T_4095_re = _RAND_7800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7801 = {1{`RANDOM}};
  _T_4095_im = _RAND_7801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7802 = {1{`RANDOM}};
  _T_4096_re = _RAND_7802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7803 = {1{`RANDOM}};
  _T_4096_im = _RAND_7803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7804 = {1{`RANDOM}};
  _T_4097_re = _RAND_7804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7805 = {1{`RANDOM}};
  _T_4097_im = _RAND_7805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7806 = {1{`RANDOM}};
  _T_4098_re = _RAND_7806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7807 = {1{`RANDOM}};
  _T_4098_im = _RAND_7807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7808 = {1{`RANDOM}};
  _T_4099_re = _RAND_7808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7809 = {1{`RANDOM}};
  _T_4099_im = _RAND_7809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7810 = {1{`RANDOM}};
  _T_4100_re = _RAND_7810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7811 = {1{`RANDOM}};
  _T_4100_im = _RAND_7811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7812 = {1{`RANDOM}};
  _T_4101_re = _RAND_7812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7813 = {1{`RANDOM}};
  _T_4101_im = _RAND_7813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7814 = {1{`RANDOM}};
  _T_4102_re = _RAND_7814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7815 = {1{`RANDOM}};
  _T_4102_im = _RAND_7815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7816 = {1{`RANDOM}};
  _T_4103_re = _RAND_7816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7817 = {1{`RANDOM}};
  _T_4103_im = _RAND_7817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7818 = {1{`RANDOM}};
  _T_4104_re = _RAND_7818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7819 = {1{`RANDOM}};
  _T_4104_im = _RAND_7819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7820 = {1{`RANDOM}};
  _T_4105_re = _RAND_7820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7821 = {1{`RANDOM}};
  _T_4105_im = _RAND_7821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7822 = {1{`RANDOM}};
  _T_4106_re = _RAND_7822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7823 = {1{`RANDOM}};
  _T_4106_im = _RAND_7823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7824 = {1{`RANDOM}};
  _T_4107_re = _RAND_7824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7825 = {1{`RANDOM}};
  _T_4107_im = _RAND_7825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7826 = {1{`RANDOM}};
  _T_4108_re = _RAND_7826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7827 = {1{`RANDOM}};
  _T_4108_im = _RAND_7827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7828 = {1{`RANDOM}};
  _T_4109_re = _RAND_7828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7829 = {1{`RANDOM}};
  _T_4109_im = _RAND_7829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7830 = {1{`RANDOM}};
  _T_4110_re = _RAND_7830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7831 = {1{`RANDOM}};
  _T_4110_im = _RAND_7831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7832 = {1{`RANDOM}};
  _T_4111_re = _RAND_7832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7833 = {1{`RANDOM}};
  _T_4111_im = _RAND_7833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7834 = {1{`RANDOM}};
  _T_4112_re = _RAND_7834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7835 = {1{`RANDOM}};
  _T_4112_im = _RAND_7835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7836 = {1{`RANDOM}};
  _T_4113_re = _RAND_7836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7837 = {1{`RANDOM}};
  _T_4113_im = _RAND_7837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7838 = {1{`RANDOM}};
  _T_4114_re = _RAND_7838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7839 = {1{`RANDOM}};
  _T_4114_im = _RAND_7839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7840 = {1{`RANDOM}};
  _T_4115_re = _RAND_7840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7841 = {1{`RANDOM}};
  _T_4115_im = _RAND_7841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7842 = {1{`RANDOM}};
  _T_4116_re = _RAND_7842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7843 = {1{`RANDOM}};
  _T_4116_im = _RAND_7843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7844 = {1{`RANDOM}};
  _T_4117_re = _RAND_7844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7845 = {1{`RANDOM}};
  _T_4117_im = _RAND_7845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7846 = {1{`RANDOM}};
  _T_4118_re = _RAND_7846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7847 = {1{`RANDOM}};
  _T_4118_im = _RAND_7847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7848 = {1{`RANDOM}};
  _T_4119_re = _RAND_7848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7849 = {1{`RANDOM}};
  _T_4119_im = _RAND_7849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7850 = {1{`RANDOM}};
  _T_4120_re = _RAND_7850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7851 = {1{`RANDOM}};
  _T_4120_im = _RAND_7851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7852 = {1{`RANDOM}};
  _T_4121_re = _RAND_7852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7853 = {1{`RANDOM}};
  _T_4121_im = _RAND_7853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7854 = {1{`RANDOM}};
  _T_4122_re = _RAND_7854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7855 = {1{`RANDOM}};
  _T_4122_im = _RAND_7855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7856 = {1{`RANDOM}};
  _T_4123_re = _RAND_7856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7857 = {1{`RANDOM}};
  _T_4123_im = _RAND_7857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7858 = {1{`RANDOM}};
  _T_4124_re = _RAND_7858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7859 = {1{`RANDOM}};
  _T_4124_im = _RAND_7859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7860 = {1{`RANDOM}};
  _T_4125_re = _RAND_7860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7861 = {1{`RANDOM}};
  _T_4125_im = _RAND_7861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7862 = {1{`RANDOM}};
  _T_4126_re = _RAND_7862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7863 = {1{`RANDOM}};
  _T_4126_im = _RAND_7863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7864 = {1{`RANDOM}};
  _T_4127_re = _RAND_7864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7865 = {1{`RANDOM}};
  _T_4127_im = _RAND_7865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7866 = {1{`RANDOM}};
  _T_4128_re = _RAND_7866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7867 = {1{`RANDOM}};
  _T_4128_im = _RAND_7867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7868 = {1{`RANDOM}};
  _T_4129_re = _RAND_7868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7869 = {1{`RANDOM}};
  _T_4129_im = _RAND_7869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7870 = {1{`RANDOM}};
  _T_4130_re = _RAND_7870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7871 = {1{`RANDOM}};
  _T_4130_im = _RAND_7871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7872 = {1{`RANDOM}};
  _T_4131_re = _RAND_7872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7873 = {1{`RANDOM}};
  _T_4131_im = _RAND_7873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7874 = {1{`RANDOM}};
  _T_4132_re = _RAND_7874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7875 = {1{`RANDOM}};
  _T_4132_im = _RAND_7875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7876 = {1{`RANDOM}};
  _T_4133_re = _RAND_7876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7877 = {1{`RANDOM}};
  _T_4133_im = _RAND_7877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7878 = {1{`RANDOM}};
  _T_4134_re = _RAND_7878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7879 = {1{`RANDOM}};
  _T_4134_im = _RAND_7879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7880 = {1{`RANDOM}};
  _T_4135_re = _RAND_7880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7881 = {1{`RANDOM}};
  _T_4135_im = _RAND_7881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7882 = {1{`RANDOM}};
  _T_4136_re = _RAND_7882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7883 = {1{`RANDOM}};
  _T_4136_im = _RAND_7883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7884 = {1{`RANDOM}};
  _T_4137_re = _RAND_7884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7885 = {1{`RANDOM}};
  _T_4137_im = _RAND_7885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7886 = {1{`RANDOM}};
  _T_4138_re = _RAND_7886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7887 = {1{`RANDOM}};
  _T_4138_im = _RAND_7887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7888 = {1{`RANDOM}};
  _T_4139_re = _RAND_7888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7889 = {1{`RANDOM}};
  _T_4139_im = _RAND_7889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7890 = {1{`RANDOM}};
  _T_4140_re = _RAND_7890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7891 = {1{`RANDOM}};
  _T_4140_im = _RAND_7891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7892 = {1{`RANDOM}};
  _T_4141_re = _RAND_7892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7893 = {1{`RANDOM}};
  _T_4141_im = _RAND_7893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7894 = {1{`RANDOM}};
  _T_4142_re = _RAND_7894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7895 = {1{`RANDOM}};
  _T_4142_im = _RAND_7895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7896 = {1{`RANDOM}};
  _T_4143_re = _RAND_7896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7897 = {1{`RANDOM}};
  _T_4143_im = _RAND_7897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7898 = {1{`RANDOM}};
  _T_4144_re = _RAND_7898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7899 = {1{`RANDOM}};
  _T_4144_im = _RAND_7899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7900 = {1{`RANDOM}};
  _T_4145_re = _RAND_7900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7901 = {1{`RANDOM}};
  _T_4145_im = _RAND_7901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7902 = {1{`RANDOM}};
  _T_4146_re = _RAND_7902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7903 = {1{`RANDOM}};
  _T_4146_im = _RAND_7903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7904 = {1{`RANDOM}};
  _T_4147_re = _RAND_7904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7905 = {1{`RANDOM}};
  _T_4147_im = _RAND_7905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7906 = {1{`RANDOM}};
  _T_4148_re = _RAND_7906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7907 = {1{`RANDOM}};
  _T_4148_im = _RAND_7907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7908 = {1{`RANDOM}};
  _T_4149_re = _RAND_7908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7909 = {1{`RANDOM}};
  _T_4149_im = _RAND_7909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7910 = {1{`RANDOM}};
  _T_4150_re = _RAND_7910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7911 = {1{`RANDOM}};
  _T_4150_im = _RAND_7911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7912 = {1{`RANDOM}};
  _T_4151_re = _RAND_7912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7913 = {1{`RANDOM}};
  _T_4151_im = _RAND_7913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7914 = {1{`RANDOM}};
  _T_4152_re = _RAND_7914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7915 = {1{`RANDOM}};
  _T_4152_im = _RAND_7915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7916 = {1{`RANDOM}};
  _T_4153_re = _RAND_7916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7917 = {1{`RANDOM}};
  _T_4153_im = _RAND_7917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7918 = {1{`RANDOM}};
  _T_4154_re = _RAND_7918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7919 = {1{`RANDOM}};
  _T_4154_im = _RAND_7919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7920 = {1{`RANDOM}};
  _T_4155_re = _RAND_7920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7921 = {1{`RANDOM}};
  _T_4155_im = _RAND_7921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7922 = {1{`RANDOM}};
  _T_4156_re = _RAND_7922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7923 = {1{`RANDOM}};
  _T_4156_im = _RAND_7923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7924 = {1{`RANDOM}};
  _T_4157_re = _RAND_7924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7925 = {1{`RANDOM}};
  _T_4157_im = _RAND_7925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7926 = {1{`RANDOM}};
  _T_4158_re = _RAND_7926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7927 = {1{`RANDOM}};
  _T_4158_im = _RAND_7927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7928 = {1{`RANDOM}};
  _T_4159_re = _RAND_7928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7929 = {1{`RANDOM}};
  _T_4159_im = _RAND_7929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7930 = {1{`RANDOM}};
  _T_4160_re = _RAND_7930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7931 = {1{`RANDOM}};
  _T_4160_im = _RAND_7931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7932 = {1{`RANDOM}};
  _T_4161_re = _RAND_7932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7933 = {1{`RANDOM}};
  _T_4161_im = _RAND_7933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7934 = {1{`RANDOM}};
  _T_4162_re = _RAND_7934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7935 = {1{`RANDOM}};
  _T_4162_im = _RAND_7935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7936 = {1{`RANDOM}};
  _T_4163_re = _RAND_7936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7937 = {1{`RANDOM}};
  _T_4163_im = _RAND_7937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7938 = {1{`RANDOM}};
  _T_4164_re = _RAND_7938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7939 = {1{`RANDOM}};
  _T_4164_im = _RAND_7939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7940 = {1{`RANDOM}};
  _T_4165_re = _RAND_7940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7941 = {1{`RANDOM}};
  _T_4165_im = _RAND_7941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7942 = {1{`RANDOM}};
  _T_4166_re = _RAND_7942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7943 = {1{`RANDOM}};
  _T_4166_im = _RAND_7943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7944 = {1{`RANDOM}};
  _T_4167_re = _RAND_7944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7945 = {1{`RANDOM}};
  _T_4167_im = _RAND_7945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7946 = {1{`RANDOM}};
  _T_4168_re = _RAND_7946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7947 = {1{`RANDOM}};
  _T_4168_im = _RAND_7947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7948 = {1{`RANDOM}};
  _T_4169_re = _RAND_7948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7949 = {1{`RANDOM}};
  _T_4169_im = _RAND_7949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7950 = {1{`RANDOM}};
  _T_4170_re = _RAND_7950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7951 = {1{`RANDOM}};
  _T_4170_im = _RAND_7951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7952 = {1{`RANDOM}};
  _T_4171_re = _RAND_7952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7953 = {1{`RANDOM}};
  _T_4171_im = _RAND_7953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7954 = {1{`RANDOM}};
  _T_4172_re = _RAND_7954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7955 = {1{`RANDOM}};
  _T_4172_im = _RAND_7955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7956 = {1{`RANDOM}};
  _T_4173_re = _RAND_7956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7957 = {1{`RANDOM}};
  _T_4173_im = _RAND_7957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7958 = {1{`RANDOM}};
  _T_4174_re = _RAND_7958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7959 = {1{`RANDOM}};
  _T_4174_im = _RAND_7959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7960 = {1{`RANDOM}};
  _T_4175_re = _RAND_7960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7961 = {1{`RANDOM}};
  _T_4175_im = _RAND_7961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7962 = {1{`RANDOM}};
  _T_4176_re = _RAND_7962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7963 = {1{`RANDOM}};
  _T_4176_im = _RAND_7963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7964 = {1{`RANDOM}};
  _T_4177_re = _RAND_7964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7965 = {1{`RANDOM}};
  _T_4177_im = _RAND_7965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7966 = {1{`RANDOM}};
  _T_4178_re = _RAND_7966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7967 = {1{`RANDOM}};
  _T_4178_im = _RAND_7967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7968 = {1{`RANDOM}};
  _T_4179_re = _RAND_7968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7969 = {1{`RANDOM}};
  _T_4179_im = _RAND_7969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7970 = {1{`RANDOM}};
  _T_4180_re = _RAND_7970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7971 = {1{`RANDOM}};
  _T_4180_im = _RAND_7971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7972 = {1{`RANDOM}};
  _T_4181_re = _RAND_7972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7973 = {1{`RANDOM}};
  _T_4181_im = _RAND_7973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7974 = {1{`RANDOM}};
  _T_4182_re = _RAND_7974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7975 = {1{`RANDOM}};
  _T_4182_im = _RAND_7975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7976 = {1{`RANDOM}};
  _T_4183_re = _RAND_7976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7977 = {1{`RANDOM}};
  _T_4183_im = _RAND_7977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7978 = {1{`RANDOM}};
  _T_4184_re = _RAND_7978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7979 = {1{`RANDOM}};
  _T_4184_im = _RAND_7979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7980 = {1{`RANDOM}};
  _T_4185_re = _RAND_7980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7981 = {1{`RANDOM}};
  _T_4185_im = _RAND_7981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7982 = {1{`RANDOM}};
  _T_4186_re = _RAND_7982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7983 = {1{`RANDOM}};
  _T_4186_im = _RAND_7983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7984 = {1{`RANDOM}};
  _T_4187_re = _RAND_7984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7985 = {1{`RANDOM}};
  _T_4187_im = _RAND_7985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7986 = {1{`RANDOM}};
  _T_4188_re = _RAND_7986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7987 = {1{`RANDOM}};
  _T_4188_im = _RAND_7987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7988 = {1{`RANDOM}};
  _T_4189_re = _RAND_7988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7989 = {1{`RANDOM}};
  _T_4189_im = _RAND_7989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7990 = {1{`RANDOM}};
  _T_4190_re = _RAND_7990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7991 = {1{`RANDOM}};
  _T_4190_im = _RAND_7991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7992 = {1{`RANDOM}};
  _T_4191_re = _RAND_7992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7993 = {1{`RANDOM}};
  _T_4191_im = _RAND_7993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7994 = {1{`RANDOM}};
  _T_4192_re = _RAND_7994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7995 = {1{`RANDOM}};
  _T_4192_im = _RAND_7995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7996 = {1{`RANDOM}};
  _T_4193_re = _RAND_7996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7997 = {1{`RANDOM}};
  _T_4193_im = _RAND_7997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7998 = {1{`RANDOM}};
  _T_4194_re = _RAND_7998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7999 = {1{`RANDOM}};
  _T_4194_im = _RAND_7999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8000 = {1{`RANDOM}};
  _T_4195_re = _RAND_8000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8001 = {1{`RANDOM}};
  _T_4195_im = _RAND_8001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8002 = {1{`RANDOM}};
  _T_4196_re = _RAND_8002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8003 = {1{`RANDOM}};
  _T_4196_im = _RAND_8003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8004 = {1{`RANDOM}};
  _T_4197_re = _RAND_8004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8005 = {1{`RANDOM}};
  _T_4197_im = _RAND_8005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8006 = {1{`RANDOM}};
  _T_4198_re = _RAND_8006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8007 = {1{`RANDOM}};
  _T_4198_im = _RAND_8007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8008 = {1{`RANDOM}};
  _T_4199_re = _RAND_8008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8009 = {1{`RANDOM}};
  _T_4199_im = _RAND_8009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8010 = {1{`RANDOM}};
  _T_4200_re = _RAND_8010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8011 = {1{`RANDOM}};
  _T_4200_im = _RAND_8011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8012 = {1{`RANDOM}};
  _T_4201_re = _RAND_8012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8013 = {1{`RANDOM}};
  _T_4201_im = _RAND_8013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8014 = {1{`RANDOM}};
  _T_4202_re = _RAND_8014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8015 = {1{`RANDOM}};
  _T_4202_im = _RAND_8015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8016 = {1{`RANDOM}};
  _T_4203_re = _RAND_8016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8017 = {1{`RANDOM}};
  _T_4203_im = _RAND_8017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8018 = {1{`RANDOM}};
  _T_4204_re = _RAND_8018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8019 = {1{`RANDOM}};
  _T_4204_im = _RAND_8019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8020 = {1{`RANDOM}};
  _T_4205_re = _RAND_8020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8021 = {1{`RANDOM}};
  _T_4205_im = _RAND_8021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8022 = {1{`RANDOM}};
  _T_4206_re = _RAND_8022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8023 = {1{`RANDOM}};
  _T_4206_im = _RAND_8023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8024 = {1{`RANDOM}};
  _T_4207_re = _RAND_8024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8025 = {1{`RANDOM}};
  _T_4207_im = _RAND_8025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8026 = {1{`RANDOM}};
  _T_4208_re = _RAND_8026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8027 = {1{`RANDOM}};
  _T_4208_im = _RAND_8027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8028 = {1{`RANDOM}};
  _T_4209_re = _RAND_8028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8029 = {1{`RANDOM}};
  _T_4209_im = _RAND_8029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8030 = {1{`RANDOM}};
  _T_4210_re = _RAND_8030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8031 = {1{`RANDOM}};
  _T_4210_im = _RAND_8031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8032 = {1{`RANDOM}};
  _T_4211_re = _RAND_8032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8033 = {1{`RANDOM}};
  _T_4211_im = _RAND_8033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8034 = {1{`RANDOM}};
  _T_4212_re = _RAND_8034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8035 = {1{`RANDOM}};
  _T_4212_im = _RAND_8035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8036 = {1{`RANDOM}};
  _T_4213_re = _RAND_8036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8037 = {1{`RANDOM}};
  _T_4213_im = _RAND_8037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8038 = {1{`RANDOM}};
  _T_4214_re = _RAND_8038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8039 = {1{`RANDOM}};
  _T_4214_im = _RAND_8039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8040 = {1{`RANDOM}};
  _T_4215_re = _RAND_8040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8041 = {1{`RANDOM}};
  _T_4215_im = _RAND_8041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8042 = {1{`RANDOM}};
  _T_4216_re = _RAND_8042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8043 = {1{`RANDOM}};
  _T_4216_im = _RAND_8043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8044 = {1{`RANDOM}};
  _T_4217_re = _RAND_8044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8045 = {1{`RANDOM}};
  _T_4217_im = _RAND_8045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8046 = {1{`RANDOM}};
  _T_4218_re = _RAND_8046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8047 = {1{`RANDOM}};
  _T_4218_im = _RAND_8047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8048 = {1{`RANDOM}};
  _T_4219_re = _RAND_8048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8049 = {1{`RANDOM}};
  _T_4219_im = _RAND_8049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8050 = {1{`RANDOM}};
  _T_4220_re = _RAND_8050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8051 = {1{`RANDOM}};
  _T_4220_im = _RAND_8051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8052 = {1{`RANDOM}};
  _T_4221_re = _RAND_8052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8053 = {1{`RANDOM}};
  _T_4221_im = _RAND_8053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8054 = {1{`RANDOM}};
  _T_4222_re = _RAND_8054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8055 = {1{`RANDOM}};
  _T_4222_im = _RAND_8055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8056 = {1{`RANDOM}};
  _T_4223_re = _RAND_8056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8057 = {1{`RANDOM}};
  _T_4223_im = _RAND_8057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8058 = {1{`RANDOM}};
  _T_4224_re = _RAND_8058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8059 = {1{`RANDOM}};
  _T_4224_im = _RAND_8059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8060 = {1{`RANDOM}};
  _T_4225_re = _RAND_8060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8061 = {1{`RANDOM}};
  _T_4225_im = _RAND_8061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8062 = {1{`RANDOM}};
  _T_4226_re = _RAND_8062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8063 = {1{`RANDOM}};
  _T_4226_im = _RAND_8063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8064 = {1{`RANDOM}};
  _T_4227_re = _RAND_8064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8065 = {1{`RANDOM}};
  _T_4227_im = _RAND_8065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8066 = {1{`RANDOM}};
  _T_4228_re = _RAND_8066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8067 = {1{`RANDOM}};
  _T_4228_im = _RAND_8067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8068 = {1{`RANDOM}};
  _T_4229_re = _RAND_8068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8069 = {1{`RANDOM}};
  _T_4229_im = _RAND_8069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8070 = {1{`RANDOM}};
  _T_4230_re = _RAND_8070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8071 = {1{`RANDOM}};
  _T_4230_im = _RAND_8071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8072 = {1{`RANDOM}};
  _T_4231_re = _RAND_8072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8073 = {1{`RANDOM}};
  _T_4231_im = _RAND_8073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8074 = {1{`RANDOM}};
  _T_4232_re = _RAND_8074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8075 = {1{`RANDOM}};
  _T_4232_im = _RAND_8075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8076 = {1{`RANDOM}};
  _T_4233_re = _RAND_8076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8077 = {1{`RANDOM}};
  _T_4233_im = _RAND_8077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8078 = {1{`RANDOM}};
  _T_4234_re = _RAND_8078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8079 = {1{`RANDOM}};
  _T_4234_im = _RAND_8079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8080 = {1{`RANDOM}};
  _T_4235_re = _RAND_8080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8081 = {1{`RANDOM}};
  _T_4235_im = _RAND_8081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8082 = {1{`RANDOM}};
  _T_4236_re = _RAND_8082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8083 = {1{`RANDOM}};
  _T_4236_im = _RAND_8083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8084 = {1{`RANDOM}};
  _T_4237_re = _RAND_8084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8085 = {1{`RANDOM}};
  _T_4237_im = _RAND_8085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8086 = {1{`RANDOM}};
  _T_4238_re = _RAND_8086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8087 = {1{`RANDOM}};
  _T_4238_im = _RAND_8087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8088 = {1{`RANDOM}};
  _T_4239_re = _RAND_8088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8089 = {1{`RANDOM}};
  _T_4239_im = _RAND_8089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8090 = {1{`RANDOM}};
  _T_4240_re = _RAND_8090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8091 = {1{`RANDOM}};
  _T_4240_im = _RAND_8091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8092 = {1{`RANDOM}};
  _T_4241_re = _RAND_8092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8093 = {1{`RANDOM}};
  _T_4241_im = _RAND_8093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8094 = {1{`RANDOM}};
  _T_4242_re = _RAND_8094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8095 = {1{`RANDOM}};
  _T_4242_im = _RAND_8095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8096 = {1{`RANDOM}};
  _T_4243_re = _RAND_8096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8097 = {1{`RANDOM}};
  _T_4243_im = _RAND_8097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8098 = {1{`RANDOM}};
  _T_4244_re = _RAND_8098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8099 = {1{`RANDOM}};
  _T_4244_im = _RAND_8099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8100 = {1{`RANDOM}};
  _T_4245_re = _RAND_8100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8101 = {1{`RANDOM}};
  _T_4245_im = _RAND_8101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8102 = {1{`RANDOM}};
  _T_4246_re = _RAND_8102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8103 = {1{`RANDOM}};
  _T_4246_im = _RAND_8103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8104 = {1{`RANDOM}};
  _T_4247_re = _RAND_8104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8105 = {1{`RANDOM}};
  _T_4247_im = _RAND_8105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8106 = {1{`RANDOM}};
  _T_4248_re = _RAND_8106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8107 = {1{`RANDOM}};
  _T_4248_im = _RAND_8107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8108 = {1{`RANDOM}};
  _T_4249_re = _RAND_8108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8109 = {1{`RANDOM}};
  _T_4249_im = _RAND_8109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8110 = {1{`RANDOM}};
  _T_4250_re = _RAND_8110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8111 = {1{`RANDOM}};
  _T_4250_im = _RAND_8111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8112 = {1{`RANDOM}};
  _T_4251_re = _RAND_8112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8113 = {1{`RANDOM}};
  _T_4251_im = _RAND_8113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8114 = {1{`RANDOM}};
  _T_4252_re = _RAND_8114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8115 = {1{`RANDOM}};
  _T_4252_im = _RAND_8115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8116 = {1{`RANDOM}};
  _T_4253_re = _RAND_8116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8117 = {1{`RANDOM}};
  _T_4253_im = _RAND_8117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8118 = {1{`RANDOM}};
  _T_4254_re = _RAND_8118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8119 = {1{`RANDOM}};
  _T_4254_im = _RAND_8119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8120 = {1{`RANDOM}};
  _T_4255_re = _RAND_8120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8121 = {1{`RANDOM}};
  _T_4255_im = _RAND_8121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8122 = {1{`RANDOM}};
  _T_4256_re = _RAND_8122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8123 = {1{`RANDOM}};
  _T_4256_im = _RAND_8123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8124 = {1{`RANDOM}};
  _T_4257_re = _RAND_8124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8125 = {1{`RANDOM}};
  _T_4257_im = _RAND_8125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8126 = {1{`RANDOM}};
  _T_4258_re = _RAND_8126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8127 = {1{`RANDOM}};
  _T_4258_im = _RAND_8127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8128 = {1{`RANDOM}};
  _T_4259_re = _RAND_8128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8129 = {1{`RANDOM}};
  _T_4259_im = _RAND_8129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8130 = {1{`RANDOM}};
  _T_4260_re = _RAND_8130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8131 = {1{`RANDOM}};
  _T_4260_im = _RAND_8131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8132 = {1{`RANDOM}};
  _T_4261_re = _RAND_8132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8133 = {1{`RANDOM}};
  _T_4261_im = _RAND_8133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8134 = {1{`RANDOM}};
  _T_4262_re = _RAND_8134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8135 = {1{`RANDOM}};
  _T_4262_im = _RAND_8135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8136 = {1{`RANDOM}};
  _T_4263_re = _RAND_8136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8137 = {1{`RANDOM}};
  _T_4263_im = _RAND_8137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8138 = {1{`RANDOM}};
  _T_4264_re = _RAND_8138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8139 = {1{`RANDOM}};
  _T_4264_im = _RAND_8139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8140 = {1{`RANDOM}};
  _T_4265_re = _RAND_8140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8141 = {1{`RANDOM}};
  _T_4265_im = _RAND_8141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8142 = {1{`RANDOM}};
  _T_4266_re = _RAND_8142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8143 = {1{`RANDOM}};
  _T_4266_im = _RAND_8143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8144 = {1{`RANDOM}};
  _T_4267_re = _RAND_8144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8145 = {1{`RANDOM}};
  _T_4267_im = _RAND_8145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8146 = {1{`RANDOM}};
  _T_4268_re = _RAND_8146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8147 = {1{`RANDOM}};
  _T_4268_im = _RAND_8147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8148 = {1{`RANDOM}};
  _T_4269_re = _RAND_8148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8149 = {1{`RANDOM}};
  _T_4269_im = _RAND_8149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8150 = {1{`RANDOM}};
  _T_4270_re = _RAND_8150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8151 = {1{`RANDOM}};
  _T_4270_im = _RAND_8151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8152 = {1{`RANDOM}};
  _T_4271_re = _RAND_8152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8153 = {1{`RANDOM}};
  _T_4271_im = _RAND_8153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8154 = {1{`RANDOM}};
  _T_4272_re = _RAND_8154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8155 = {1{`RANDOM}};
  _T_4272_im = _RAND_8155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8156 = {1{`RANDOM}};
  _T_4273_re = _RAND_8156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8157 = {1{`RANDOM}};
  _T_4273_im = _RAND_8157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8158 = {1{`RANDOM}};
  _T_4274_re = _RAND_8158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8159 = {1{`RANDOM}};
  _T_4274_im = _RAND_8159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8160 = {1{`RANDOM}};
  _T_4275_re = _RAND_8160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8161 = {1{`RANDOM}};
  _T_4275_im = _RAND_8161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8162 = {1{`RANDOM}};
  _T_4276_re = _RAND_8162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8163 = {1{`RANDOM}};
  _T_4276_im = _RAND_8163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8164 = {1{`RANDOM}};
  _T_4277_re = _RAND_8164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8165 = {1{`RANDOM}};
  _T_4277_im = _RAND_8165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8166 = {1{`RANDOM}};
  _T_4278_re = _RAND_8166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8167 = {1{`RANDOM}};
  _T_4278_im = _RAND_8167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8168 = {1{`RANDOM}};
  _T_4279_re = _RAND_8168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8169 = {1{`RANDOM}};
  _T_4279_im = _RAND_8169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8170 = {1{`RANDOM}};
  _T_4280_re = _RAND_8170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8171 = {1{`RANDOM}};
  _T_4280_im = _RAND_8171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8172 = {1{`RANDOM}};
  _T_4281_re = _RAND_8172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8173 = {1{`RANDOM}};
  _T_4281_im = _RAND_8173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8174 = {1{`RANDOM}};
  _T_4282_re = _RAND_8174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8175 = {1{`RANDOM}};
  _T_4282_im = _RAND_8175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8176 = {1{`RANDOM}};
  _T_4283_re = _RAND_8176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8177 = {1{`RANDOM}};
  _T_4283_im = _RAND_8177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8178 = {1{`RANDOM}};
  _T_4284_re = _RAND_8178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8179 = {1{`RANDOM}};
  _T_4284_im = _RAND_8179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8180 = {1{`RANDOM}};
  _T_4285_re = _RAND_8180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8181 = {1{`RANDOM}};
  _T_4285_im = _RAND_8181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8182 = {1{`RANDOM}};
  _T_4286_re = _RAND_8182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8183 = {1{`RANDOM}};
  _T_4286_im = _RAND_8183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8184 = {1{`RANDOM}};
  _T_4287_re = _RAND_8184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8185 = {1{`RANDOM}};
  _T_4287_im = _RAND_8185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8186 = {1{`RANDOM}};
  _T_4288_re = _RAND_8186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8187 = {1{`RANDOM}};
  _T_4288_im = _RAND_8187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8188 = {1{`RANDOM}};
  _T_4289_re = _RAND_8188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8189 = {1{`RANDOM}};
  _T_4289_im = _RAND_8189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8190 = {1{`RANDOM}};
  _T_4290_re = _RAND_8190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8191 = {1{`RANDOM}};
  _T_4290_im = _RAND_8191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8192 = {1{`RANDOM}};
  _T_4291_re = _RAND_8192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8193 = {1{`RANDOM}};
  _T_4291_im = _RAND_8193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8194 = {1{`RANDOM}};
  _T_4294_re = _RAND_8194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8195 = {1{`RANDOM}};
  _T_4294_im = _RAND_8195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8196 = {1{`RANDOM}};
  _T_4295_re = _RAND_8196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8197 = {1{`RANDOM}};
  _T_4295_im = _RAND_8197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8198 = {1{`RANDOM}};
  _T_4296_re = _RAND_8198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8199 = {1{`RANDOM}};
  _T_4296_im = _RAND_8199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8200 = {1{`RANDOM}};
  _T_4297_re = _RAND_8200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8201 = {1{`RANDOM}};
  _T_4297_im = _RAND_8201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8202 = {1{`RANDOM}};
  _T_4298_re = _RAND_8202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8203 = {1{`RANDOM}};
  _T_4298_im = _RAND_8203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8204 = {1{`RANDOM}};
  _T_4299_re = _RAND_8204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8205 = {1{`RANDOM}};
  _T_4299_im = _RAND_8205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8206 = {1{`RANDOM}};
  _T_4300_re = _RAND_8206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8207 = {1{`RANDOM}};
  _T_4300_im = _RAND_8207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8208 = {1{`RANDOM}};
  _T_4301_re = _RAND_8208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8209 = {1{`RANDOM}};
  _T_4301_im = _RAND_8209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8210 = {1{`RANDOM}};
  _T_4302_re = _RAND_8210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8211 = {1{`RANDOM}};
  _T_4302_im = _RAND_8211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8212 = {1{`RANDOM}};
  _T_4303_re = _RAND_8212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8213 = {1{`RANDOM}};
  _T_4303_im = _RAND_8213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8214 = {1{`RANDOM}};
  _T_4304_re = _RAND_8214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8215 = {1{`RANDOM}};
  _T_4304_im = _RAND_8215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8216 = {1{`RANDOM}};
  _T_4305_re = _RAND_8216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8217 = {1{`RANDOM}};
  _T_4305_im = _RAND_8217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8218 = {1{`RANDOM}};
  _T_4306_re = _RAND_8218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8219 = {1{`RANDOM}};
  _T_4306_im = _RAND_8219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8220 = {1{`RANDOM}};
  _T_4307_re = _RAND_8220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8221 = {1{`RANDOM}};
  _T_4307_im = _RAND_8221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8222 = {1{`RANDOM}};
  _T_4308_re = _RAND_8222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8223 = {1{`RANDOM}};
  _T_4308_im = _RAND_8223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8224 = {1{`RANDOM}};
  _T_4309_re = _RAND_8224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8225 = {1{`RANDOM}};
  _T_4309_im = _RAND_8225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8226 = {1{`RANDOM}};
  _T_4310_re = _RAND_8226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8227 = {1{`RANDOM}};
  _T_4310_im = _RAND_8227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8228 = {1{`RANDOM}};
  _T_4311_re = _RAND_8228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8229 = {1{`RANDOM}};
  _T_4311_im = _RAND_8229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8230 = {1{`RANDOM}};
  _T_4312_re = _RAND_8230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8231 = {1{`RANDOM}};
  _T_4312_im = _RAND_8231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8232 = {1{`RANDOM}};
  _T_4313_re = _RAND_8232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8233 = {1{`RANDOM}};
  _T_4313_im = _RAND_8233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8234 = {1{`RANDOM}};
  _T_4314_re = _RAND_8234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8235 = {1{`RANDOM}};
  _T_4314_im = _RAND_8235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8236 = {1{`RANDOM}};
  _T_4315_re = _RAND_8236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8237 = {1{`RANDOM}};
  _T_4315_im = _RAND_8237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8238 = {1{`RANDOM}};
  _T_4316_re = _RAND_8238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8239 = {1{`RANDOM}};
  _T_4316_im = _RAND_8239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8240 = {1{`RANDOM}};
  _T_4317_re = _RAND_8240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8241 = {1{`RANDOM}};
  _T_4317_im = _RAND_8241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8242 = {1{`RANDOM}};
  _T_4318_re = _RAND_8242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8243 = {1{`RANDOM}};
  _T_4318_im = _RAND_8243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8244 = {1{`RANDOM}};
  _T_4319_re = _RAND_8244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8245 = {1{`RANDOM}};
  _T_4319_im = _RAND_8245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8246 = {1{`RANDOM}};
  _T_4320_re = _RAND_8246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8247 = {1{`RANDOM}};
  _T_4320_im = _RAND_8247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8248 = {1{`RANDOM}};
  _T_4321_re = _RAND_8248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8249 = {1{`RANDOM}};
  _T_4321_im = _RAND_8249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8250 = {1{`RANDOM}};
  _T_4322_re = _RAND_8250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8251 = {1{`RANDOM}};
  _T_4322_im = _RAND_8251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8252 = {1{`RANDOM}};
  _T_4323_re = _RAND_8252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8253 = {1{`RANDOM}};
  _T_4323_im = _RAND_8253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8254 = {1{`RANDOM}};
  _T_4324_re = _RAND_8254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8255 = {1{`RANDOM}};
  _T_4324_im = _RAND_8255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8256 = {1{`RANDOM}};
  _T_4325_re = _RAND_8256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8257 = {1{`RANDOM}};
  _T_4325_im = _RAND_8257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8258 = {1{`RANDOM}};
  _T_4326_re = _RAND_8258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8259 = {1{`RANDOM}};
  _T_4326_im = _RAND_8259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8260 = {1{`RANDOM}};
  _T_4327_re = _RAND_8260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8261 = {1{`RANDOM}};
  _T_4327_im = _RAND_8261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8262 = {1{`RANDOM}};
  _T_4328_re = _RAND_8262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8263 = {1{`RANDOM}};
  _T_4328_im = _RAND_8263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8264 = {1{`RANDOM}};
  _T_4329_re = _RAND_8264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8265 = {1{`RANDOM}};
  _T_4329_im = _RAND_8265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8266 = {1{`RANDOM}};
  _T_4330_re = _RAND_8266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8267 = {1{`RANDOM}};
  _T_4330_im = _RAND_8267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8268 = {1{`RANDOM}};
  _T_4331_re = _RAND_8268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8269 = {1{`RANDOM}};
  _T_4331_im = _RAND_8269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8270 = {1{`RANDOM}};
  _T_4332_re = _RAND_8270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8271 = {1{`RANDOM}};
  _T_4332_im = _RAND_8271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8272 = {1{`RANDOM}};
  _T_4333_re = _RAND_8272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8273 = {1{`RANDOM}};
  _T_4333_im = _RAND_8273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8274 = {1{`RANDOM}};
  _T_4334_re = _RAND_8274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8275 = {1{`RANDOM}};
  _T_4334_im = _RAND_8275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8276 = {1{`RANDOM}};
  _T_4335_re = _RAND_8276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8277 = {1{`RANDOM}};
  _T_4335_im = _RAND_8277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8278 = {1{`RANDOM}};
  _T_4336_re = _RAND_8278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8279 = {1{`RANDOM}};
  _T_4336_im = _RAND_8279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8280 = {1{`RANDOM}};
  _T_4337_re = _RAND_8280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8281 = {1{`RANDOM}};
  _T_4337_im = _RAND_8281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8282 = {1{`RANDOM}};
  _T_4338_re = _RAND_8282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8283 = {1{`RANDOM}};
  _T_4338_im = _RAND_8283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8284 = {1{`RANDOM}};
  _T_4339_re = _RAND_8284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8285 = {1{`RANDOM}};
  _T_4339_im = _RAND_8285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8286 = {1{`RANDOM}};
  _T_4340_re = _RAND_8286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8287 = {1{`RANDOM}};
  _T_4340_im = _RAND_8287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8288 = {1{`RANDOM}};
  _T_4341_re = _RAND_8288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8289 = {1{`RANDOM}};
  _T_4341_im = _RAND_8289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8290 = {1{`RANDOM}};
  _T_4342_re = _RAND_8290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8291 = {1{`RANDOM}};
  _T_4342_im = _RAND_8291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8292 = {1{`RANDOM}};
  _T_4343_re = _RAND_8292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8293 = {1{`RANDOM}};
  _T_4343_im = _RAND_8293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8294 = {1{`RANDOM}};
  _T_4344_re = _RAND_8294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8295 = {1{`RANDOM}};
  _T_4344_im = _RAND_8295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8296 = {1{`RANDOM}};
  _T_4345_re = _RAND_8296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8297 = {1{`RANDOM}};
  _T_4345_im = _RAND_8297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8298 = {1{`RANDOM}};
  _T_4346_re = _RAND_8298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8299 = {1{`RANDOM}};
  _T_4346_im = _RAND_8299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8300 = {1{`RANDOM}};
  _T_4347_re = _RAND_8300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8301 = {1{`RANDOM}};
  _T_4347_im = _RAND_8301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8302 = {1{`RANDOM}};
  _T_4348_re = _RAND_8302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8303 = {1{`RANDOM}};
  _T_4348_im = _RAND_8303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8304 = {1{`RANDOM}};
  _T_4349_re = _RAND_8304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8305 = {1{`RANDOM}};
  _T_4349_im = _RAND_8305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8306 = {1{`RANDOM}};
  _T_4350_re = _RAND_8306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8307 = {1{`RANDOM}};
  _T_4350_im = _RAND_8307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8308 = {1{`RANDOM}};
  _T_4351_re = _RAND_8308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8309 = {1{`RANDOM}};
  _T_4351_im = _RAND_8309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8310 = {1{`RANDOM}};
  _T_4352_re = _RAND_8310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8311 = {1{`RANDOM}};
  _T_4352_im = _RAND_8311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8312 = {1{`RANDOM}};
  _T_4353_re = _RAND_8312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8313 = {1{`RANDOM}};
  _T_4353_im = _RAND_8313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8314 = {1{`RANDOM}};
  _T_4354_re = _RAND_8314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8315 = {1{`RANDOM}};
  _T_4354_im = _RAND_8315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8316 = {1{`RANDOM}};
  _T_4355_re = _RAND_8316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8317 = {1{`RANDOM}};
  _T_4355_im = _RAND_8317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8318 = {1{`RANDOM}};
  _T_4356_re = _RAND_8318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8319 = {1{`RANDOM}};
  _T_4356_im = _RAND_8319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8320 = {1{`RANDOM}};
  _T_4357_re = _RAND_8320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8321 = {1{`RANDOM}};
  _T_4357_im = _RAND_8321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8322 = {1{`RANDOM}};
  _T_4358_re = _RAND_8322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8323 = {1{`RANDOM}};
  _T_4358_im = _RAND_8323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8324 = {1{`RANDOM}};
  _T_4359_re = _RAND_8324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8325 = {1{`RANDOM}};
  _T_4359_im = _RAND_8325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8326 = {1{`RANDOM}};
  _T_4360_re = _RAND_8326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8327 = {1{`RANDOM}};
  _T_4360_im = _RAND_8327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8328 = {1{`RANDOM}};
  _T_4361_re = _RAND_8328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8329 = {1{`RANDOM}};
  _T_4361_im = _RAND_8329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8330 = {1{`RANDOM}};
  _T_4362_re = _RAND_8330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8331 = {1{`RANDOM}};
  _T_4362_im = _RAND_8331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8332 = {1{`RANDOM}};
  _T_4363_re = _RAND_8332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8333 = {1{`RANDOM}};
  _T_4363_im = _RAND_8333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8334 = {1{`RANDOM}};
  _T_4364_re = _RAND_8334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8335 = {1{`RANDOM}};
  _T_4364_im = _RAND_8335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8336 = {1{`RANDOM}};
  _T_4365_re = _RAND_8336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8337 = {1{`RANDOM}};
  _T_4365_im = _RAND_8337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8338 = {1{`RANDOM}};
  _T_4366_re = _RAND_8338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8339 = {1{`RANDOM}};
  _T_4366_im = _RAND_8339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8340 = {1{`RANDOM}};
  _T_4367_re = _RAND_8340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8341 = {1{`RANDOM}};
  _T_4367_im = _RAND_8341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8342 = {1{`RANDOM}};
  _T_4368_re = _RAND_8342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8343 = {1{`RANDOM}};
  _T_4368_im = _RAND_8343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8344 = {1{`RANDOM}};
  _T_4369_re = _RAND_8344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8345 = {1{`RANDOM}};
  _T_4369_im = _RAND_8345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8346 = {1{`RANDOM}};
  _T_4370_re = _RAND_8346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8347 = {1{`RANDOM}};
  _T_4370_im = _RAND_8347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8348 = {1{`RANDOM}};
  _T_4371_re = _RAND_8348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8349 = {1{`RANDOM}};
  _T_4371_im = _RAND_8349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8350 = {1{`RANDOM}};
  _T_4372_re = _RAND_8350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8351 = {1{`RANDOM}};
  _T_4372_im = _RAND_8351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8352 = {1{`RANDOM}};
  _T_4373_re = _RAND_8352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8353 = {1{`RANDOM}};
  _T_4373_im = _RAND_8353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8354 = {1{`RANDOM}};
  _T_4374_re = _RAND_8354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8355 = {1{`RANDOM}};
  _T_4374_im = _RAND_8355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8356 = {1{`RANDOM}};
  _T_4375_re = _RAND_8356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8357 = {1{`RANDOM}};
  _T_4375_im = _RAND_8357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8358 = {1{`RANDOM}};
  _T_4376_re = _RAND_8358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8359 = {1{`RANDOM}};
  _T_4376_im = _RAND_8359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8360 = {1{`RANDOM}};
  _T_4377_re = _RAND_8360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8361 = {1{`RANDOM}};
  _T_4377_im = _RAND_8361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8362 = {1{`RANDOM}};
  _T_4378_re = _RAND_8362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8363 = {1{`RANDOM}};
  _T_4378_im = _RAND_8363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8364 = {1{`RANDOM}};
  _T_4379_re = _RAND_8364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8365 = {1{`RANDOM}};
  _T_4379_im = _RAND_8365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8366 = {1{`RANDOM}};
  _T_4380_re = _RAND_8366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8367 = {1{`RANDOM}};
  _T_4380_im = _RAND_8367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8368 = {1{`RANDOM}};
  _T_4381_re = _RAND_8368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8369 = {1{`RANDOM}};
  _T_4381_im = _RAND_8369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8370 = {1{`RANDOM}};
  _T_4382_re = _RAND_8370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8371 = {1{`RANDOM}};
  _T_4382_im = _RAND_8371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8372 = {1{`RANDOM}};
  _T_4383_re = _RAND_8372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8373 = {1{`RANDOM}};
  _T_4383_im = _RAND_8373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8374 = {1{`RANDOM}};
  _T_4384_re = _RAND_8374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8375 = {1{`RANDOM}};
  _T_4384_im = _RAND_8375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8376 = {1{`RANDOM}};
  _T_4385_re = _RAND_8376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8377 = {1{`RANDOM}};
  _T_4385_im = _RAND_8377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8378 = {1{`RANDOM}};
  _T_4386_re = _RAND_8378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8379 = {1{`RANDOM}};
  _T_4386_im = _RAND_8379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8380 = {1{`RANDOM}};
  _T_4387_re = _RAND_8380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8381 = {1{`RANDOM}};
  _T_4387_im = _RAND_8381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8382 = {1{`RANDOM}};
  _T_4388_re = _RAND_8382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8383 = {1{`RANDOM}};
  _T_4388_im = _RAND_8383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8384 = {1{`RANDOM}};
  _T_4389_re = _RAND_8384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8385 = {1{`RANDOM}};
  _T_4389_im = _RAND_8385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8386 = {1{`RANDOM}};
  _T_4390_re = _RAND_8386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8387 = {1{`RANDOM}};
  _T_4390_im = _RAND_8387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8388 = {1{`RANDOM}};
  _T_4391_re = _RAND_8388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8389 = {1{`RANDOM}};
  _T_4391_im = _RAND_8389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8390 = {1{`RANDOM}};
  _T_4392_re = _RAND_8390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8391 = {1{`RANDOM}};
  _T_4392_im = _RAND_8391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8392 = {1{`RANDOM}};
  _T_4393_re = _RAND_8392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8393 = {1{`RANDOM}};
  _T_4393_im = _RAND_8393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8394 = {1{`RANDOM}};
  _T_4394_re = _RAND_8394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8395 = {1{`RANDOM}};
  _T_4394_im = _RAND_8395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8396 = {1{`RANDOM}};
  _T_4395_re = _RAND_8396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8397 = {1{`RANDOM}};
  _T_4395_im = _RAND_8397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8398 = {1{`RANDOM}};
  _T_4396_re = _RAND_8398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8399 = {1{`RANDOM}};
  _T_4396_im = _RAND_8399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8400 = {1{`RANDOM}};
  _T_4397_re = _RAND_8400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8401 = {1{`RANDOM}};
  _T_4397_im = _RAND_8401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8402 = {1{`RANDOM}};
  _T_4398_re = _RAND_8402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8403 = {1{`RANDOM}};
  _T_4398_im = _RAND_8403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8404 = {1{`RANDOM}};
  _T_4399_re = _RAND_8404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8405 = {1{`RANDOM}};
  _T_4399_im = _RAND_8405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8406 = {1{`RANDOM}};
  _T_4400_re = _RAND_8406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8407 = {1{`RANDOM}};
  _T_4400_im = _RAND_8407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8408 = {1{`RANDOM}};
  _T_4401_re = _RAND_8408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8409 = {1{`RANDOM}};
  _T_4401_im = _RAND_8409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8410 = {1{`RANDOM}};
  _T_4402_re = _RAND_8410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8411 = {1{`RANDOM}};
  _T_4402_im = _RAND_8411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8412 = {1{`RANDOM}};
  _T_4403_re = _RAND_8412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8413 = {1{`RANDOM}};
  _T_4403_im = _RAND_8413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8414 = {1{`RANDOM}};
  _T_4404_re = _RAND_8414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8415 = {1{`RANDOM}};
  _T_4404_im = _RAND_8415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8416 = {1{`RANDOM}};
  _T_4405_re = _RAND_8416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8417 = {1{`RANDOM}};
  _T_4405_im = _RAND_8417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8418 = {1{`RANDOM}};
  _T_4406_re = _RAND_8418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8419 = {1{`RANDOM}};
  _T_4406_im = _RAND_8419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8420 = {1{`RANDOM}};
  _T_4407_re = _RAND_8420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8421 = {1{`RANDOM}};
  _T_4407_im = _RAND_8421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8422 = {1{`RANDOM}};
  _T_4408_re = _RAND_8422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8423 = {1{`RANDOM}};
  _T_4408_im = _RAND_8423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8424 = {1{`RANDOM}};
  _T_4409_re = _RAND_8424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8425 = {1{`RANDOM}};
  _T_4409_im = _RAND_8425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8426 = {1{`RANDOM}};
  _T_4410_re = _RAND_8426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8427 = {1{`RANDOM}};
  _T_4410_im = _RAND_8427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8428 = {1{`RANDOM}};
  _T_4411_re = _RAND_8428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8429 = {1{`RANDOM}};
  _T_4411_im = _RAND_8429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8430 = {1{`RANDOM}};
  _T_4412_re = _RAND_8430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8431 = {1{`RANDOM}};
  _T_4412_im = _RAND_8431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8432 = {1{`RANDOM}};
  _T_4413_re = _RAND_8432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8433 = {1{`RANDOM}};
  _T_4413_im = _RAND_8433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8434 = {1{`RANDOM}};
  _T_4414_re = _RAND_8434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8435 = {1{`RANDOM}};
  _T_4414_im = _RAND_8435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8436 = {1{`RANDOM}};
  _T_4415_re = _RAND_8436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8437 = {1{`RANDOM}};
  _T_4415_im = _RAND_8437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8438 = {1{`RANDOM}};
  _T_4416_re = _RAND_8438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8439 = {1{`RANDOM}};
  _T_4416_im = _RAND_8439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8440 = {1{`RANDOM}};
  _T_4417_re = _RAND_8440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8441 = {1{`RANDOM}};
  _T_4417_im = _RAND_8441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8442 = {1{`RANDOM}};
  _T_4418_re = _RAND_8442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8443 = {1{`RANDOM}};
  _T_4418_im = _RAND_8443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8444 = {1{`RANDOM}};
  _T_4419_re = _RAND_8444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8445 = {1{`RANDOM}};
  _T_4419_im = _RAND_8445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8446 = {1{`RANDOM}};
  _T_4420_re = _RAND_8446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8447 = {1{`RANDOM}};
  _T_4420_im = _RAND_8447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8448 = {1{`RANDOM}};
  _T_4421_re = _RAND_8448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8449 = {1{`RANDOM}};
  _T_4421_im = _RAND_8449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8450 = {1{`RANDOM}};
  _T_4422_re = _RAND_8450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8451 = {1{`RANDOM}};
  _T_4422_im = _RAND_8451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8452 = {1{`RANDOM}};
  _T_4423_re = _RAND_8452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8453 = {1{`RANDOM}};
  _T_4423_im = _RAND_8453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8454 = {1{`RANDOM}};
  _T_4424_re = _RAND_8454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8455 = {1{`RANDOM}};
  _T_4424_im = _RAND_8455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8456 = {1{`RANDOM}};
  _T_4425_re = _RAND_8456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8457 = {1{`RANDOM}};
  _T_4425_im = _RAND_8457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8458 = {1{`RANDOM}};
  _T_4426_re = _RAND_8458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8459 = {1{`RANDOM}};
  _T_4426_im = _RAND_8459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8460 = {1{`RANDOM}};
  _T_4427_re = _RAND_8460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8461 = {1{`RANDOM}};
  _T_4427_im = _RAND_8461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8462 = {1{`RANDOM}};
  _T_4428_re = _RAND_8462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8463 = {1{`RANDOM}};
  _T_4428_im = _RAND_8463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8464 = {1{`RANDOM}};
  _T_4429_re = _RAND_8464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8465 = {1{`RANDOM}};
  _T_4429_im = _RAND_8465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8466 = {1{`RANDOM}};
  _T_4430_re = _RAND_8466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8467 = {1{`RANDOM}};
  _T_4430_im = _RAND_8467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8468 = {1{`RANDOM}};
  _T_4431_re = _RAND_8468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8469 = {1{`RANDOM}};
  _T_4431_im = _RAND_8469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8470 = {1{`RANDOM}};
  _T_4432_re = _RAND_8470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8471 = {1{`RANDOM}};
  _T_4432_im = _RAND_8471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8472 = {1{`RANDOM}};
  _T_4433_re = _RAND_8472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8473 = {1{`RANDOM}};
  _T_4433_im = _RAND_8473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8474 = {1{`RANDOM}};
  _T_4434_re = _RAND_8474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8475 = {1{`RANDOM}};
  _T_4434_im = _RAND_8475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8476 = {1{`RANDOM}};
  _T_4435_re = _RAND_8476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8477 = {1{`RANDOM}};
  _T_4435_im = _RAND_8477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8478 = {1{`RANDOM}};
  _T_4436_re = _RAND_8478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8479 = {1{`RANDOM}};
  _T_4436_im = _RAND_8479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8480 = {1{`RANDOM}};
  _T_4437_re = _RAND_8480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8481 = {1{`RANDOM}};
  _T_4437_im = _RAND_8481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8482 = {1{`RANDOM}};
  _T_4438_re = _RAND_8482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8483 = {1{`RANDOM}};
  _T_4438_im = _RAND_8483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8484 = {1{`RANDOM}};
  _T_4439_re = _RAND_8484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8485 = {1{`RANDOM}};
  _T_4439_im = _RAND_8485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8486 = {1{`RANDOM}};
  _T_4440_re = _RAND_8486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8487 = {1{`RANDOM}};
  _T_4440_im = _RAND_8487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8488 = {1{`RANDOM}};
  _T_4441_re = _RAND_8488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8489 = {1{`RANDOM}};
  _T_4441_im = _RAND_8489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8490 = {1{`RANDOM}};
  _T_4442_re = _RAND_8490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8491 = {1{`RANDOM}};
  _T_4442_im = _RAND_8491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8492 = {1{`RANDOM}};
  _T_4443_re = _RAND_8492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8493 = {1{`RANDOM}};
  _T_4443_im = _RAND_8493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8494 = {1{`RANDOM}};
  _T_4444_re = _RAND_8494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8495 = {1{`RANDOM}};
  _T_4444_im = _RAND_8495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8496 = {1{`RANDOM}};
  _T_4445_re = _RAND_8496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8497 = {1{`RANDOM}};
  _T_4445_im = _RAND_8497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8498 = {1{`RANDOM}};
  _T_4446_re = _RAND_8498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8499 = {1{`RANDOM}};
  _T_4446_im = _RAND_8499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8500 = {1{`RANDOM}};
  _T_4447_re = _RAND_8500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8501 = {1{`RANDOM}};
  _T_4447_im = _RAND_8501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8502 = {1{`RANDOM}};
  _T_4448_re = _RAND_8502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8503 = {1{`RANDOM}};
  _T_4448_im = _RAND_8503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8504 = {1{`RANDOM}};
  _T_4449_re = _RAND_8504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8505 = {1{`RANDOM}};
  _T_4449_im = _RAND_8505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8506 = {1{`RANDOM}};
  _T_4450_re = _RAND_8506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8507 = {1{`RANDOM}};
  _T_4450_im = _RAND_8507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8508 = {1{`RANDOM}};
  _T_4451_re = _RAND_8508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8509 = {1{`RANDOM}};
  _T_4451_im = _RAND_8509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8510 = {1{`RANDOM}};
  _T_4452_re = _RAND_8510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8511 = {1{`RANDOM}};
  _T_4452_im = _RAND_8511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8512 = {1{`RANDOM}};
  _T_4453_re = _RAND_8512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8513 = {1{`RANDOM}};
  _T_4453_im = _RAND_8513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8514 = {1{`RANDOM}};
  _T_4454_re = _RAND_8514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8515 = {1{`RANDOM}};
  _T_4454_im = _RAND_8515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8516 = {1{`RANDOM}};
  _T_4455_re = _RAND_8516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8517 = {1{`RANDOM}};
  _T_4455_im = _RAND_8517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8518 = {1{`RANDOM}};
  _T_4456_re = _RAND_8518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8519 = {1{`RANDOM}};
  _T_4456_im = _RAND_8519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8520 = {1{`RANDOM}};
  _T_4457_re = _RAND_8520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8521 = {1{`RANDOM}};
  _T_4457_im = _RAND_8521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8522 = {1{`RANDOM}};
  _T_4458_re = _RAND_8522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8523 = {1{`RANDOM}};
  _T_4458_im = _RAND_8523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8524 = {1{`RANDOM}};
  _T_4459_re = _RAND_8524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8525 = {1{`RANDOM}};
  _T_4459_im = _RAND_8525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8526 = {1{`RANDOM}};
  _T_4460_re = _RAND_8526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8527 = {1{`RANDOM}};
  _T_4460_im = _RAND_8527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8528 = {1{`RANDOM}};
  _T_4461_re = _RAND_8528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8529 = {1{`RANDOM}};
  _T_4461_im = _RAND_8529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8530 = {1{`RANDOM}};
  _T_4462_re = _RAND_8530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8531 = {1{`RANDOM}};
  _T_4462_im = _RAND_8531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8532 = {1{`RANDOM}};
  _T_4463_re = _RAND_8532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8533 = {1{`RANDOM}};
  _T_4463_im = _RAND_8533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8534 = {1{`RANDOM}};
  _T_4464_re = _RAND_8534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8535 = {1{`RANDOM}};
  _T_4464_im = _RAND_8535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8536 = {1{`RANDOM}};
  _T_4465_re = _RAND_8536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8537 = {1{`RANDOM}};
  _T_4465_im = _RAND_8537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8538 = {1{`RANDOM}};
  _T_4466_re = _RAND_8538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8539 = {1{`RANDOM}};
  _T_4466_im = _RAND_8539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8540 = {1{`RANDOM}};
  _T_4467_re = _RAND_8540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8541 = {1{`RANDOM}};
  _T_4467_im = _RAND_8541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8542 = {1{`RANDOM}};
  _T_4468_re = _RAND_8542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8543 = {1{`RANDOM}};
  _T_4468_im = _RAND_8543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8544 = {1{`RANDOM}};
  _T_4469_re = _RAND_8544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8545 = {1{`RANDOM}};
  _T_4469_im = _RAND_8545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8546 = {1{`RANDOM}};
  _T_4470_re = _RAND_8546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8547 = {1{`RANDOM}};
  _T_4470_im = _RAND_8547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8548 = {1{`RANDOM}};
  _T_4471_re = _RAND_8548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8549 = {1{`RANDOM}};
  _T_4471_im = _RAND_8549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8550 = {1{`RANDOM}};
  _T_4472_re = _RAND_8550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8551 = {1{`RANDOM}};
  _T_4472_im = _RAND_8551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8552 = {1{`RANDOM}};
  _T_4473_re = _RAND_8552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8553 = {1{`RANDOM}};
  _T_4473_im = _RAND_8553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8554 = {1{`RANDOM}};
  _T_4474_re = _RAND_8554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8555 = {1{`RANDOM}};
  _T_4474_im = _RAND_8555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8556 = {1{`RANDOM}};
  _T_4475_re = _RAND_8556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8557 = {1{`RANDOM}};
  _T_4475_im = _RAND_8557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8558 = {1{`RANDOM}};
  _T_4476_re = _RAND_8558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8559 = {1{`RANDOM}};
  _T_4476_im = _RAND_8559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8560 = {1{`RANDOM}};
  _T_4477_re = _RAND_8560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8561 = {1{`RANDOM}};
  _T_4477_im = _RAND_8561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8562 = {1{`RANDOM}};
  _T_4478_re = _RAND_8562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8563 = {1{`RANDOM}};
  _T_4478_im = _RAND_8563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8564 = {1{`RANDOM}};
  _T_4479_re = _RAND_8564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8565 = {1{`RANDOM}};
  _T_4479_im = _RAND_8565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8566 = {1{`RANDOM}};
  _T_4480_re = _RAND_8566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8567 = {1{`RANDOM}};
  _T_4480_im = _RAND_8567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8568 = {1{`RANDOM}};
  _T_4481_re = _RAND_8568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8569 = {1{`RANDOM}};
  _T_4481_im = _RAND_8569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8570 = {1{`RANDOM}};
  _T_4482_re = _RAND_8570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8571 = {1{`RANDOM}};
  _T_4482_im = _RAND_8571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8572 = {1{`RANDOM}};
  _T_4483_re = _RAND_8572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8573 = {1{`RANDOM}};
  _T_4483_im = _RAND_8573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8574 = {1{`RANDOM}};
  _T_4484_re = _RAND_8574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8575 = {1{`RANDOM}};
  _T_4484_im = _RAND_8575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8576 = {1{`RANDOM}};
  _T_4485_re = _RAND_8576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8577 = {1{`RANDOM}};
  _T_4485_im = _RAND_8577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8578 = {1{`RANDOM}};
  _T_4486_re = _RAND_8578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8579 = {1{`RANDOM}};
  _T_4486_im = _RAND_8579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8580 = {1{`RANDOM}};
  _T_4487_re = _RAND_8580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8581 = {1{`RANDOM}};
  _T_4487_im = _RAND_8581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8582 = {1{`RANDOM}};
  _T_4488_re = _RAND_8582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8583 = {1{`RANDOM}};
  _T_4488_im = _RAND_8583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8584 = {1{`RANDOM}};
  _T_4489_re = _RAND_8584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8585 = {1{`RANDOM}};
  _T_4489_im = _RAND_8585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8586 = {1{`RANDOM}};
  _T_4490_re = _RAND_8586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8587 = {1{`RANDOM}};
  _T_4490_im = _RAND_8587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8588 = {1{`RANDOM}};
  _T_4491_re = _RAND_8588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8589 = {1{`RANDOM}};
  _T_4491_im = _RAND_8589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8590 = {1{`RANDOM}};
  _T_4492_re = _RAND_8590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8591 = {1{`RANDOM}};
  _T_4492_im = _RAND_8591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8592 = {1{`RANDOM}};
  _T_4493_re = _RAND_8592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8593 = {1{`RANDOM}};
  _T_4493_im = _RAND_8593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8594 = {1{`RANDOM}};
  _T_4494_re = _RAND_8594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8595 = {1{`RANDOM}};
  _T_4494_im = _RAND_8595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8596 = {1{`RANDOM}};
  _T_4495_re = _RAND_8596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8597 = {1{`RANDOM}};
  _T_4495_im = _RAND_8597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8598 = {1{`RANDOM}};
  _T_4496_re = _RAND_8598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8599 = {1{`RANDOM}};
  _T_4496_im = _RAND_8599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8600 = {1{`RANDOM}};
  _T_4497_re = _RAND_8600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8601 = {1{`RANDOM}};
  _T_4497_im = _RAND_8601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8602 = {1{`RANDOM}};
  _T_4498_re = _RAND_8602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8603 = {1{`RANDOM}};
  _T_4498_im = _RAND_8603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8604 = {1{`RANDOM}};
  _T_4499_re = _RAND_8604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8605 = {1{`RANDOM}};
  _T_4499_im = _RAND_8605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8606 = {1{`RANDOM}};
  _T_4500_re = _RAND_8606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8607 = {1{`RANDOM}};
  _T_4500_im = _RAND_8607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8608 = {1{`RANDOM}};
  _T_4501_re = _RAND_8608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8609 = {1{`RANDOM}};
  _T_4501_im = _RAND_8609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8610 = {1{`RANDOM}};
  _T_4502_re = _RAND_8610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8611 = {1{`RANDOM}};
  _T_4502_im = _RAND_8611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8612 = {1{`RANDOM}};
  _T_4503_re = _RAND_8612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8613 = {1{`RANDOM}};
  _T_4503_im = _RAND_8613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8614 = {1{`RANDOM}};
  _T_4504_re = _RAND_8614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8615 = {1{`RANDOM}};
  _T_4504_im = _RAND_8615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8616 = {1{`RANDOM}};
  _T_4505_re = _RAND_8616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8617 = {1{`RANDOM}};
  _T_4505_im = _RAND_8617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8618 = {1{`RANDOM}};
  _T_4506_re = _RAND_8618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8619 = {1{`RANDOM}};
  _T_4506_im = _RAND_8619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8620 = {1{`RANDOM}};
  _T_4507_re = _RAND_8620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8621 = {1{`RANDOM}};
  _T_4507_im = _RAND_8621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8622 = {1{`RANDOM}};
  _T_4508_re = _RAND_8622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8623 = {1{`RANDOM}};
  _T_4508_im = _RAND_8623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8624 = {1{`RANDOM}};
  _T_4509_re = _RAND_8624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8625 = {1{`RANDOM}};
  _T_4509_im = _RAND_8625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8626 = {1{`RANDOM}};
  _T_4510_re = _RAND_8626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8627 = {1{`RANDOM}};
  _T_4510_im = _RAND_8627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8628 = {1{`RANDOM}};
  _T_4511_re = _RAND_8628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8629 = {1{`RANDOM}};
  _T_4511_im = _RAND_8629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8630 = {1{`RANDOM}};
  _T_4512_re = _RAND_8630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8631 = {1{`RANDOM}};
  _T_4512_im = _RAND_8631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8632 = {1{`RANDOM}};
  _T_4513_re = _RAND_8632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8633 = {1{`RANDOM}};
  _T_4513_im = _RAND_8633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8634 = {1{`RANDOM}};
  _T_4514_re = _RAND_8634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8635 = {1{`RANDOM}};
  _T_4514_im = _RAND_8635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8636 = {1{`RANDOM}};
  _T_4515_re = _RAND_8636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8637 = {1{`RANDOM}};
  _T_4515_im = _RAND_8637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8638 = {1{`RANDOM}};
  _T_4516_re = _RAND_8638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8639 = {1{`RANDOM}};
  _T_4516_im = _RAND_8639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8640 = {1{`RANDOM}};
  _T_4517_re = _RAND_8640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8641 = {1{`RANDOM}};
  _T_4517_im = _RAND_8641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8642 = {1{`RANDOM}};
  _T_4518_re = _RAND_8642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8643 = {1{`RANDOM}};
  _T_4518_im = _RAND_8643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8644 = {1{`RANDOM}};
  _T_4519_re = _RAND_8644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8645 = {1{`RANDOM}};
  _T_4519_im = _RAND_8645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8646 = {1{`RANDOM}};
  _T_4520_re = _RAND_8646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8647 = {1{`RANDOM}};
  _T_4520_im = _RAND_8647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8648 = {1{`RANDOM}};
  _T_4521_re = _RAND_8648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8649 = {1{`RANDOM}};
  _T_4521_im = _RAND_8649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8650 = {1{`RANDOM}};
  _T_4522_re = _RAND_8650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8651 = {1{`RANDOM}};
  _T_4522_im = _RAND_8651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8652 = {1{`RANDOM}};
  _T_4523_re = _RAND_8652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8653 = {1{`RANDOM}};
  _T_4523_im = _RAND_8653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8654 = {1{`RANDOM}};
  _T_4524_re = _RAND_8654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8655 = {1{`RANDOM}};
  _T_4524_im = _RAND_8655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8656 = {1{`RANDOM}};
  _T_4525_re = _RAND_8656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8657 = {1{`RANDOM}};
  _T_4525_im = _RAND_8657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8658 = {1{`RANDOM}};
  _T_4526_re = _RAND_8658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8659 = {1{`RANDOM}};
  _T_4526_im = _RAND_8659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8660 = {1{`RANDOM}};
  _T_4527_re = _RAND_8660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8661 = {1{`RANDOM}};
  _T_4527_im = _RAND_8661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8662 = {1{`RANDOM}};
  _T_4528_re = _RAND_8662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8663 = {1{`RANDOM}};
  _T_4528_im = _RAND_8663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8664 = {1{`RANDOM}};
  _T_4529_re = _RAND_8664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8665 = {1{`RANDOM}};
  _T_4529_im = _RAND_8665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8666 = {1{`RANDOM}};
  _T_4530_re = _RAND_8666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8667 = {1{`RANDOM}};
  _T_4530_im = _RAND_8667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8668 = {1{`RANDOM}};
  _T_4531_re = _RAND_8668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8669 = {1{`RANDOM}};
  _T_4531_im = _RAND_8669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8670 = {1{`RANDOM}};
  _T_4532_re = _RAND_8670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8671 = {1{`RANDOM}};
  _T_4532_im = _RAND_8671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8672 = {1{`RANDOM}};
  _T_4533_re = _RAND_8672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8673 = {1{`RANDOM}};
  _T_4533_im = _RAND_8673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8674 = {1{`RANDOM}};
  _T_4534_re = _RAND_8674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8675 = {1{`RANDOM}};
  _T_4534_im = _RAND_8675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8676 = {1{`RANDOM}};
  _T_4535_re = _RAND_8676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8677 = {1{`RANDOM}};
  _T_4535_im = _RAND_8677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8678 = {1{`RANDOM}};
  _T_4536_re = _RAND_8678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8679 = {1{`RANDOM}};
  _T_4536_im = _RAND_8679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8680 = {1{`RANDOM}};
  _T_4537_re = _RAND_8680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8681 = {1{`RANDOM}};
  _T_4537_im = _RAND_8681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8682 = {1{`RANDOM}};
  _T_4538_re = _RAND_8682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8683 = {1{`RANDOM}};
  _T_4538_im = _RAND_8683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8684 = {1{`RANDOM}};
  _T_4539_re = _RAND_8684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8685 = {1{`RANDOM}};
  _T_4539_im = _RAND_8685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8686 = {1{`RANDOM}};
  _T_4540_re = _RAND_8686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8687 = {1{`RANDOM}};
  _T_4540_im = _RAND_8687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8688 = {1{`RANDOM}};
  _T_4541_re = _RAND_8688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8689 = {1{`RANDOM}};
  _T_4541_im = _RAND_8689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8690 = {1{`RANDOM}};
  _T_4542_re = _RAND_8690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8691 = {1{`RANDOM}};
  _T_4542_im = _RAND_8691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8692 = {1{`RANDOM}};
  _T_4543_re = _RAND_8692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8693 = {1{`RANDOM}};
  _T_4543_im = _RAND_8693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8694 = {1{`RANDOM}};
  _T_4544_re = _RAND_8694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8695 = {1{`RANDOM}};
  _T_4544_im = _RAND_8695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8696 = {1{`RANDOM}};
  _T_4545_re = _RAND_8696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8697 = {1{`RANDOM}};
  _T_4545_im = _RAND_8697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8698 = {1{`RANDOM}};
  _T_4546_re = _RAND_8698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8699 = {1{`RANDOM}};
  _T_4546_im = _RAND_8699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8700 = {1{`RANDOM}};
  _T_4547_re = _RAND_8700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8701 = {1{`RANDOM}};
  _T_4547_im = _RAND_8701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8702 = {1{`RANDOM}};
  _T_4548_re = _RAND_8702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8703 = {1{`RANDOM}};
  _T_4548_im = _RAND_8703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8704 = {1{`RANDOM}};
  _T_4549_re = _RAND_8704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8705 = {1{`RANDOM}};
  _T_4549_im = _RAND_8705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8706 = {1{`RANDOM}};
  _T_4550_re = _RAND_8706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8707 = {1{`RANDOM}};
  _T_4550_im = _RAND_8707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8708 = {1{`RANDOM}};
  _T_4551_re = _RAND_8708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8709 = {1{`RANDOM}};
  _T_4551_im = _RAND_8709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8710 = {1{`RANDOM}};
  _T_4552_re = _RAND_8710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8711 = {1{`RANDOM}};
  _T_4552_im = _RAND_8711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8712 = {1{`RANDOM}};
  _T_4553_re = _RAND_8712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8713 = {1{`RANDOM}};
  _T_4553_im = _RAND_8713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8714 = {1{`RANDOM}};
  _T_4554_re = _RAND_8714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8715 = {1{`RANDOM}};
  _T_4554_im = _RAND_8715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8716 = {1{`RANDOM}};
  _T_4555_re = _RAND_8716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8717 = {1{`RANDOM}};
  _T_4555_im = _RAND_8717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8718 = {1{`RANDOM}};
  _T_4556_re = _RAND_8718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8719 = {1{`RANDOM}};
  _T_4556_im = _RAND_8719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8720 = {1{`RANDOM}};
  _T_4557_re = _RAND_8720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8721 = {1{`RANDOM}};
  _T_4557_im = _RAND_8721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8722 = {1{`RANDOM}};
  _T_4558_re = _RAND_8722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8723 = {1{`RANDOM}};
  _T_4558_im = _RAND_8723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8724 = {1{`RANDOM}};
  _T_4559_re = _RAND_8724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8725 = {1{`RANDOM}};
  _T_4559_im = _RAND_8725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8726 = {1{`RANDOM}};
  _T_4560_re = _RAND_8726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8727 = {1{`RANDOM}};
  _T_4560_im = _RAND_8727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8728 = {1{`RANDOM}};
  _T_4561_re = _RAND_8728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8729 = {1{`RANDOM}};
  _T_4561_im = _RAND_8729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8730 = {1{`RANDOM}};
  _T_4562_re = _RAND_8730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8731 = {1{`RANDOM}};
  _T_4562_im = _RAND_8731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8732 = {1{`RANDOM}};
  _T_4563_re = _RAND_8732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8733 = {1{`RANDOM}};
  _T_4563_im = _RAND_8733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8734 = {1{`RANDOM}};
  _T_4564_re = _RAND_8734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8735 = {1{`RANDOM}};
  _T_4564_im = _RAND_8735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8736 = {1{`RANDOM}};
  _T_4565_re = _RAND_8736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8737 = {1{`RANDOM}};
  _T_4565_im = _RAND_8737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8738 = {1{`RANDOM}};
  _T_4566_re = _RAND_8738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8739 = {1{`RANDOM}};
  _T_4566_im = _RAND_8739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8740 = {1{`RANDOM}};
  _T_4567_re = _RAND_8740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8741 = {1{`RANDOM}};
  _T_4567_im = _RAND_8741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8742 = {1{`RANDOM}};
  _T_4568_re = _RAND_8742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8743 = {1{`RANDOM}};
  _T_4568_im = _RAND_8743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8744 = {1{`RANDOM}};
  _T_4569_re = _RAND_8744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8745 = {1{`RANDOM}};
  _T_4569_im = _RAND_8745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8746 = {1{`RANDOM}};
  _T_4570_re = _RAND_8746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8747 = {1{`RANDOM}};
  _T_4570_im = _RAND_8747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8748 = {1{`RANDOM}};
  _T_4571_re = _RAND_8748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8749 = {1{`RANDOM}};
  _T_4571_im = _RAND_8749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8750 = {1{`RANDOM}};
  _T_4572_re = _RAND_8750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8751 = {1{`RANDOM}};
  _T_4572_im = _RAND_8751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8752 = {1{`RANDOM}};
  _T_4573_re = _RAND_8752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8753 = {1{`RANDOM}};
  _T_4573_im = _RAND_8753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8754 = {1{`RANDOM}};
  _T_4574_re = _RAND_8754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8755 = {1{`RANDOM}};
  _T_4574_im = _RAND_8755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8756 = {1{`RANDOM}};
  _T_4575_re = _RAND_8756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8757 = {1{`RANDOM}};
  _T_4575_im = _RAND_8757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8758 = {1{`RANDOM}};
  _T_4576_re = _RAND_8758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8759 = {1{`RANDOM}};
  _T_4576_im = _RAND_8759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8760 = {1{`RANDOM}};
  _T_4577_re = _RAND_8760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8761 = {1{`RANDOM}};
  _T_4577_im = _RAND_8761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8762 = {1{`RANDOM}};
  _T_4578_re = _RAND_8762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8763 = {1{`RANDOM}};
  _T_4578_im = _RAND_8763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8764 = {1{`RANDOM}};
  _T_4579_re = _RAND_8764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8765 = {1{`RANDOM}};
  _T_4579_im = _RAND_8765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8766 = {1{`RANDOM}};
  _T_4580_re = _RAND_8766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8767 = {1{`RANDOM}};
  _T_4580_im = _RAND_8767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8768 = {1{`RANDOM}};
  _T_4581_re = _RAND_8768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8769 = {1{`RANDOM}};
  _T_4581_im = _RAND_8769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8770 = {1{`RANDOM}};
  _T_4582_re = _RAND_8770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8771 = {1{`RANDOM}};
  _T_4582_im = _RAND_8771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8772 = {1{`RANDOM}};
  _T_4583_re = _RAND_8772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8773 = {1{`RANDOM}};
  _T_4583_im = _RAND_8773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8774 = {1{`RANDOM}};
  _T_4584_re = _RAND_8774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8775 = {1{`RANDOM}};
  _T_4584_im = _RAND_8775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8776 = {1{`RANDOM}};
  _T_4585_re = _RAND_8776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8777 = {1{`RANDOM}};
  _T_4585_im = _RAND_8777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8778 = {1{`RANDOM}};
  _T_4586_re = _RAND_8778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8779 = {1{`RANDOM}};
  _T_4586_im = _RAND_8779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8780 = {1{`RANDOM}};
  _T_4587_re = _RAND_8780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8781 = {1{`RANDOM}};
  _T_4587_im = _RAND_8781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8782 = {1{`RANDOM}};
  _T_4588_re = _RAND_8782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8783 = {1{`RANDOM}};
  _T_4588_im = _RAND_8783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8784 = {1{`RANDOM}};
  _T_4589_re = _RAND_8784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8785 = {1{`RANDOM}};
  _T_4589_im = _RAND_8785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8786 = {1{`RANDOM}};
  _T_4590_re = _RAND_8786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8787 = {1{`RANDOM}};
  _T_4590_im = _RAND_8787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8788 = {1{`RANDOM}};
  _T_4591_re = _RAND_8788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8789 = {1{`RANDOM}};
  _T_4591_im = _RAND_8789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8790 = {1{`RANDOM}};
  _T_4592_re = _RAND_8790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8791 = {1{`RANDOM}};
  _T_4592_im = _RAND_8791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8792 = {1{`RANDOM}};
  _T_4593_re = _RAND_8792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8793 = {1{`RANDOM}};
  _T_4593_im = _RAND_8793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8794 = {1{`RANDOM}};
  _T_4594_re = _RAND_8794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8795 = {1{`RANDOM}};
  _T_4594_im = _RAND_8795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8796 = {1{`RANDOM}};
  _T_4595_re = _RAND_8796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8797 = {1{`RANDOM}};
  _T_4595_im = _RAND_8797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8798 = {1{`RANDOM}};
  _T_4596_re = _RAND_8798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8799 = {1{`RANDOM}};
  _T_4596_im = _RAND_8799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8800 = {1{`RANDOM}};
  _T_4597_re = _RAND_8800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8801 = {1{`RANDOM}};
  _T_4597_im = _RAND_8801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8802 = {1{`RANDOM}};
  _T_4598_re = _RAND_8802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8803 = {1{`RANDOM}};
  _T_4598_im = _RAND_8803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8804 = {1{`RANDOM}};
  _T_4599_re = _RAND_8804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8805 = {1{`RANDOM}};
  _T_4599_im = _RAND_8805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8806 = {1{`RANDOM}};
  _T_4600_re = _RAND_8806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8807 = {1{`RANDOM}};
  _T_4600_im = _RAND_8807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8808 = {1{`RANDOM}};
  _T_4601_re = _RAND_8808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8809 = {1{`RANDOM}};
  _T_4601_im = _RAND_8809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8810 = {1{`RANDOM}};
  _T_4602_re = _RAND_8810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8811 = {1{`RANDOM}};
  _T_4602_im = _RAND_8811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8812 = {1{`RANDOM}};
  _T_4603_re = _RAND_8812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8813 = {1{`RANDOM}};
  _T_4603_im = _RAND_8813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8814 = {1{`RANDOM}};
  _T_4604_re = _RAND_8814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8815 = {1{`RANDOM}};
  _T_4604_im = _RAND_8815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8816 = {1{`RANDOM}};
  _T_4605_re = _RAND_8816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8817 = {1{`RANDOM}};
  _T_4605_im = _RAND_8817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8818 = {1{`RANDOM}};
  _T_4606_re = _RAND_8818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8819 = {1{`RANDOM}};
  _T_4606_im = _RAND_8819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8820 = {1{`RANDOM}};
  _T_4607_re = _RAND_8820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8821 = {1{`RANDOM}};
  _T_4607_im = _RAND_8821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8822 = {1{`RANDOM}};
  _T_4608_re = _RAND_8822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8823 = {1{`RANDOM}};
  _T_4608_im = _RAND_8823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8824 = {1{`RANDOM}};
  _T_4609_re = _RAND_8824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8825 = {1{`RANDOM}};
  _T_4609_im = _RAND_8825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8826 = {1{`RANDOM}};
  _T_4610_re = _RAND_8826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8827 = {1{`RANDOM}};
  _T_4610_im = _RAND_8827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8828 = {1{`RANDOM}};
  _T_4611_re = _RAND_8828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8829 = {1{`RANDOM}};
  _T_4611_im = _RAND_8829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8830 = {1{`RANDOM}};
  _T_4612_re = _RAND_8830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8831 = {1{`RANDOM}};
  _T_4612_im = _RAND_8831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8832 = {1{`RANDOM}};
  _T_4613_re = _RAND_8832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8833 = {1{`RANDOM}};
  _T_4613_im = _RAND_8833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8834 = {1{`RANDOM}};
  _T_4614_re = _RAND_8834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8835 = {1{`RANDOM}};
  _T_4614_im = _RAND_8835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8836 = {1{`RANDOM}};
  _T_4615_re = _RAND_8836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8837 = {1{`RANDOM}};
  _T_4615_im = _RAND_8837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8838 = {1{`RANDOM}};
  _T_4616_re = _RAND_8838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8839 = {1{`RANDOM}};
  _T_4616_im = _RAND_8839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8840 = {1{`RANDOM}};
  _T_4617_re = _RAND_8840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8841 = {1{`RANDOM}};
  _T_4617_im = _RAND_8841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8842 = {1{`RANDOM}};
  _T_4618_re = _RAND_8842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8843 = {1{`RANDOM}};
  _T_4618_im = _RAND_8843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8844 = {1{`RANDOM}};
  _T_4619_re = _RAND_8844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8845 = {1{`RANDOM}};
  _T_4619_im = _RAND_8845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8846 = {1{`RANDOM}};
  _T_4620_re = _RAND_8846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8847 = {1{`RANDOM}};
  _T_4620_im = _RAND_8847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8848 = {1{`RANDOM}};
  _T_4621_re = _RAND_8848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8849 = {1{`RANDOM}};
  _T_4621_im = _RAND_8849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8850 = {1{`RANDOM}};
  _T_4622_re = _RAND_8850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8851 = {1{`RANDOM}};
  _T_4622_im = _RAND_8851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8852 = {1{`RANDOM}};
  _T_4623_re = _RAND_8852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8853 = {1{`RANDOM}};
  _T_4623_im = _RAND_8853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8854 = {1{`RANDOM}};
  _T_4624_re = _RAND_8854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8855 = {1{`RANDOM}};
  _T_4624_im = _RAND_8855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8856 = {1{`RANDOM}};
  _T_4625_re = _RAND_8856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8857 = {1{`RANDOM}};
  _T_4625_im = _RAND_8857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8858 = {1{`RANDOM}};
  _T_4626_re = _RAND_8858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8859 = {1{`RANDOM}};
  _T_4626_im = _RAND_8859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8860 = {1{`RANDOM}};
  _T_4627_re = _RAND_8860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8861 = {1{`RANDOM}};
  _T_4627_im = _RAND_8861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8862 = {1{`RANDOM}};
  _T_4628_re = _RAND_8862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8863 = {1{`RANDOM}};
  _T_4628_im = _RAND_8863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8864 = {1{`RANDOM}};
  _T_4629_re = _RAND_8864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8865 = {1{`RANDOM}};
  _T_4629_im = _RAND_8865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8866 = {1{`RANDOM}};
  _T_4630_re = _RAND_8866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8867 = {1{`RANDOM}};
  _T_4630_im = _RAND_8867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8868 = {1{`RANDOM}};
  _T_4631_re = _RAND_8868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8869 = {1{`RANDOM}};
  _T_4631_im = _RAND_8869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8870 = {1{`RANDOM}};
  _T_4632_re = _RAND_8870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8871 = {1{`RANDOM}};
  _T_4632_im = _RAND_8871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8872 = {1{`RANDOM}};
  _T_4633_re = _RAND_8872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8873 = {1{`RANDOM}};
  _T_4633_im = _RAND_8873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8874 = {1{`RANDOM}};
  _T_4634_re = _RAND_8874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8875 = {1{`RANDOM}};
  _T_4634_im = _RAND_8875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8876 = {1{`RANDOM}};
  _T_4635_re = _RAND_8876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8877 = {1{`RANDOM}};
  _T_4635_im = _RAND_8877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8878 = {1{`RANDOM}};
  _T_4636_re = _RAND_8878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8879 = {1{`RANDOM}};
  _T_4636_im = _RAND_8879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8880 = {1{`RANDOM}};
  _T_4637_re = _RAND_8880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8881 = {1{`RANDOM}};
  _T_4637_im = _RAND_8881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8882 = {1{`RANDOM}};
  _T_4638_re = _RAND_8882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8883 = {1{`RANDOM}};
  _T_4638_im = _RAND_8883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8884 = {1{`RANDOM}};
  _T_4639_re = _RAND_8884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8885 = {1{`RANDOM}};
  _T_4639_im = _RAND_8885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8886 = {1{`RANDOM}};
  _T_4640_re = _RAND_8886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8887 = {1{`RANDOM}};
  _T_4640_im = _RAND_8887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8888 = {1{`RANDOM}};
  _T_4641_re = _RAND_8888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8889 = {1{`RANDOM}};
  _T_4641_im = _RAND_8889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8890 = {1{`RANDOM}};
  _T_4642_re = _RAND_8890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8891 = {1{`RANDOM}};
  _T_4642_im = _RAND_8891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8892 = {1{`RANDOM}};
  _T_4643_re = _RAND_8892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8893 = {1{`RANDOM}};
  _T_4643_im = _RAND_8893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8894 = {1{`RANDOM}};
  _T_4644_re = _RAND_8894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8895 = {1{`RANDOM}};
  _T_4644_im = _RAND_8895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8896 = {1{`RANDOM}};
  _T_4645_re = _RAND_8896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8897 = {1{`RANDOM}};
  _T_4645_im = _RAND_8897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8898 = {1{`RANDOM}};
  _T_4646_re = _RAND_8898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8899 = {1{`RANDOM}};
  _T_4646_im = _RAND_8899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8900 = {1{`RANDOM}};
  _T_4647_re = _RAND_8900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8901 = {1{`RANDOM}};
  _T_4647_im = _RAND_8901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8902 = {1{`RANDOM}};
  _T_4648_re = _RAND_8902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8903 = {1{`RANDOM}};
  _T_4648_im = _RAND_8903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8904 = {1{`RANDOM}};
  _T_4649_re = _RAND_8904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8905 = {1{`RANDOM}};
  _T_4649_im = _RAND_8905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8906 = {1{`RANDOM}};
  _T_4650_re = _RAND_8906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8907 = {1{`RANDOM}};
  _T_4650_im = _RAND_8907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8908 = {1{`RANDOM}};
  _T_4651_re = _RAND_8908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8909 = {1{`RANDOM}};
  _T_4651_im = _RAND_8909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8910 = {1{`RANDOM}};
  _T_4652_re = _RAND_8910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8911 = {1{`RANDOM}};
  _T_4652_im = _RAND_8911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8912 = {1{`RANDOM}};
  _T_4653_re = _RAND_8912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8913 = {1{`RANDOM}};
  _T_4653_im = _RAND_8913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8914 = {1{`RANDOM}};
  _T_4654_re = _RAND_8914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8915 = {1{`RANDOM}};
  _T_4654_im = _RAND_8915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8916 = {1{`RANDOM}};
  _T_4655_re = _RAND_8916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8917 = {1{`RANDOM}};
  _T_4655_im = _RAND_8917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8918 = {1{`RANDOM}};
  _T_4656_re = _RAND_8918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8919 = {1{`RANDOM}};
  _T_4656_im = _RAND_8919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8920 = {1{`RANDOM}};
  _T_4657_re = _RAND_8920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8921 = {1{`RANDOM}};
  _T_4657_im = _RAND_8921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8922 = {1{`RANDOM}};
  _T_4658_re = _RAND_8922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8923 = {1{`RANDOM}};
  _T_4658_im = _RAND_8923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8924 = {1{`RANDOM}};
  _T_4659_re = _RAND_8924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8925 = {1{`RANDOM}};
  _T_4659_im = _RAND_8925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8926 = {1{`RANDOM}};
  _T_4660_re = _RAND_8926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8927 = {1{`RANDOM}};
  _T_4660_im = _RAND_8927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8928 = {1{`RANDOM}};
  _T_4661_re = _RAND_8928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8929 = {1{`RANDOM}};
  _T_4661_im = _RAND_8929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8930 = {1{`RANDOM}};
  _T_4662_re = _RAND_8930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8931 = {1{`RANDOM}};
  _T_4662_im = _RAND_8931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8932 = {1{`RANDOM}};
  _T_4663_re = _RAND_8932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8933 = {1{`RANDOM}};
  _T_4663_im = _RAND_8933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8934 = {1{`RANDOM}};
  _T_4664_re = _RAND_8934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8935 = {1{`RANDOM}};
  _T_4664_im = _RAND_8935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8936 = {1{`RANDOM}};
  _T_4665_re = _RAND_8936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8937 = {1{`RANDOM}};
  _T_4665_im = _RAND_8937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8938 = {1{`RANDOM}};
  _T_4666_re = _RAND_8938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8939 = {1{`RANDOM}};
  _T_4666_im = _RAND_8939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8940 = {1{`RANDOM}};
  _T_4667_re = _RAND_8940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8941 = {1{`RANDOM}};
  _T_4667_im = _RAND_8941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8942 = {1{`RANDOM}};
  _T_4668_re = _RAND_8942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8943 = {1{`RANDOM}};
  _T_4668_im = _RAND_8943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8944 = {1{`RANDOM}};
  _T_4669_re = _RAND_8944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8945 = {1{`RANDOM}};
  _T_4669_im = _RAND_8945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8946 = {1{`RANDOM}};
  _T_4670_re = _RAND_8946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8947 = {1{`RANDOM}};
  _T_4670_im = _RAND_8947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8948 = {1{`RANDOM}};
  _T_4671_re = _RAND_8948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8949 = {1{`RANDOM}};
  _T_4671_im = _RAND_8949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8950 = {1{`RANDOM}};
  _T_4672_re = _RAND_8950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8951 = {1{`RANDOM}};
  _T_4672_im = _RAND_8951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8952 = {1{`RANDOM}};
  _T_4673_re = _RAND_8952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8953 = {1{`RANDOM}};
  _T_4673_im = _RAND_8953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8954 = {1{`RANDOM}};
  _T_4674_re = _RAND_8954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8955 = {1{`RANDOM}};
  _T_4674_im = _RAND_8955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8956 = {1{`RANDOM}};
  _T_4675_re = _RAND_8956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8957 = {1{`RANDOM}};
  _T_4675_im = _RAND_8957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8958 = {1{`RANDOM}};
  _T_4676_re = _RAND_8958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8959 = {1{`RANDOM}};
  _T_4676_im = _RAND_8959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8960 = {1{`RANDOM}};
  _T_4677_re = _RAND_8960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8961 = {1{`RANDOM}};
  _T_4677_im = _RAND_8961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8962 = {1{`RANDOM}};
  _T_4678_re = _RAND_8962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8963 = {1{`RANDOM}};
  _T_4678_im = _RAND_8963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8964 = {1{`RANDOM}};
  _T_4679_re = _RAND_8964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8965 = {1{`RANDOM}};
  _T_4679_im = _RAND_8965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8966 = {1{`RANDOM}};
  _T_4680_re = _RAND_8966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8967 = {1{`RANDOM}};
  _T_4680_im = _RAND_8967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8968 = {1{`RANDOM}};
  _T_4681_re = _RAND_8968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8969 = {1{`RANDOM}};
  _T_4681_im = _RAND_8969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8970 = {1{`RANDOM}};
  _T_4682_re = _RAND_8970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8971 = {1{`RANDOM}};
  _T_4682_im = _RAND_8971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8972 = {1{`RANDOM}};
  _T_4683_re = _RAND_8972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8973 = {1{`RANDOM}};
  _T_4683_im = _RAND_8973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8974 = {1{`RANDOM}};
  _T_4684_re = _RAND_8974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8975 = {1{`RANDOM}};
  _T_4684_im = _RAND_8975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8976 = {1{`RANDOM}};
  _T_4685_re = _RAND_8976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8977 = {1{`RANDOM}};
  _T_4685_im = _RAND_8977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8978 = {1{`RANDOM}};
  _T_4686_re = _RAND_8978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8979 = {1{`RANDOM}};
  _T_4686_im = _RAND_8979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8980 = {1{`RANDOM}};
  _T_4687_re = _RAND_8980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8981 = {1{`RANDOM}};
  _T_4687_im = _RAND_8981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8982 = {1{`RANDOM}};
  _T_4688_re = _RAND_8982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8983 = {1{`RANDOM}};
  _T_4688_im = _RAND_8983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8984 = {1{`RANDOM}};
  _T_4689_re = _RAND_8984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8985 = {1{`RANDOM}};
  _T_4689_im = _RAND_8985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8986 = {1{`RANDOM}};
  _T_4690_re = _RAND_8986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8987 = {1{`RANDOM}};
  _T_4690_im = _RAND_8987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8988 = {1{`RANDOM}};
  _T_4691_re = _RAND_8988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8989 = {1{`RANDOM}};
  _T_4691_im = _RAND_8989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8990 = {1{`RANDOM}};
  _T_4692_re = _RAND_8990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8991 = {1{`RANDOM}};
  _T_4692_im = _RAND_8991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8992 = {1{`RANDOM}};
  _T_4693_re = _RAND_8992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8993 = {1{`RANDOM}};
  _T_4693_im = _RAND_8993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8994 = {1{`RANDOM}};
  _T_4694_re = _RAND_8994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8995 = {1{`RANDOM}};
  _T_4694_im = _RAND_8995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8996 = {1{`RANDOM}};
  _T_4695_re = _RAND_8996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8997 = {1{`RANDOM}};
  _T_4695_im = _RAND_8997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8998 = {1{`RANDOM}};
  _T_4696_re = _RAND_8998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8999 = {1{`RANDOM}};
  _T_4696_im = _RAND_8999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9000 = {1{`RANDOM}};
  _T_4697_re = _RAND_9000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9001 = {1{`RANDOM}};
  _T_4697_im = _RAND_9001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9002 = {1{`RANDOM}};
  _T_4698_re = _RAND_9002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9003 = {1{`RANDOM}};
  _T_4698_im = _RAND_9003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9004 = {1{`RANDOM}};
  _T_4699_re = _RAND_9004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9005 = {1{`RANDOM}};
  _T_4699_im = _RAND_9005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9006 = {1{`RANDOM}};
  _T_4700_re = _RAND_9006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9007 = {1{`RANDOM}};
  _T_4700_im = _RAND_9007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9008 = {1{`RANDOM}};
  _T_4701_re = _RAND_9008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9009 = {1{`RANDOM}};
  _T_4701_im = _RAND_9009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9010 = {1{`RANDOM}};
  _T_4702_re = _RAND_9010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9011 = {1{`RANDOM}};
  _T_4702_im = _RAND_9011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9012 = {1{`RANDOM}};
  _T_4703_re = _RAND_9012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9013 = {1{`RANDOM}};
  _T_4703_im = _RAND_9013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9014 = {1{`RANDOM}};
  _T_4704_re = _RAND_9014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9015 = {1{`RANDOM}};
  _T_4704_im = _RAND_9015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9016 = {1{`RANDOM}};
  _T_4705_re = _RAND_9016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9017 = {1{`RANDOM}};
  _T_4705_im = _RAND_9017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9018 = {1{`RANDOM}};
  _T_4706_re = _RAND_9018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9019 = {1{`RANDOM}};
  _T_4706_im = _RAND_9019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9020 = {1{`RANDOM}};
  _T_4707_re = _RAND_9020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9021 = {1{`RANDOM}};
  _T_4707_im = _RAND_9021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9022 = {1{`RANDOM}};
  _T_4708_re = _RAND_9022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9023 = {1{`RANDOM}};
  _T_4708_im = _RAND_9023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9024 = {1{`RANDOM}};
  _T_4709_re = _RAND_9024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9025 = {1{`RANDOM}};
  _T_4709_im = _RAND_9025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9026 = {1{`RANDOM}};
  _T_4710_re = _RAND_9026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9027 = {1{`RANDOM}};
  _T_4710_im = _RAND_9027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9028 = {1{`RANDOM}};
  _T_4711_re = _RAND_9028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9029 = {1{`RANDOM}};
  _T_4711_im = _RAND_9029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9030 = {1{`RANDOM}};
  _T_4712_re = _RAND_9030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9031 = {1{`RANDOM}};
  _T_4712_im = _RAND_9031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9032 = {1{`RANDOM}};
  _T_4713_re = _RAND_9032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9033 = {1{`RANDOM}};
  _T_4713_im = _RAND_9033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9034 = {1{`RANDOM}};
  _T_4714_re = _RAND_9034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9035 = {1{`RANDOM}};
  _T_4714_im = _RAND_9035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9036 = {1{`RANDOM}};
  _T_4715_re = _RAND_9036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9037 = {1{`RANDOM}};
  _T_4715_im = _RAND_9037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9038 = {1{`RANDOM}};
  _T_4716_re = _RAND_9038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9039 = {1{`RANDOM}};
  _T_4716_im = _RAND_9039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9040 = {1{`RANDOM}};
  _T_4717_re = _RAND_9040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9041 = {1{`RANDOM}};
  _T_4717_im = _RAND_9041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9042 = {1{`RANDOM}};
  _T_4718_re = _RAND_9042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9043 = {1{`RANDOM}};
  _T_4718_im = _RAND_9043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9044 = {1{`RANDOM}};
  _T_4719_re = _RAND_9044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9045 = {1{`RANDOM}};
  _T_4719_im = _RAND_9045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9046 = {1{`RANDOM}};
  _T_4720_re = _RAND_9046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9047 = {1{`RANDOM}};
  _T_4720_im = _RAND_9047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9048 = {1{`RANDOM}};
  _T_4721_re = _RAND_9048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9049 = {1{`RANDOM}};
  _T_4721_im = _RAND_9049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9050 = {1{`RANDOM}};
  _T_4722_re = _RAND_9050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9051 = {1{`RANDOM}};
  _T_4722_im = _RAND_9051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9052 = {1{`RANDOM}};
  _T_4723_re = _RAND_9052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9053 = {1{`RANDOM}};
  _T_4723_im = _RAND_9053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9054 = {1{`RANDOM}};
  _T_4724_re = _RAND_9054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9055 = {1{`RANDOM}};
  _T_4724_im = _RAND_9055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9056 = {1{`RANDOM}};
  _T_4725_re = _RAND_9056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9057 = {1{`RANDOM}};
  _T_4725_im = _RAND_9057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9058 = {1{`RANDOM}};
  _T_4726_re = _RAND_9058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9059 = {1{`RANDOM}};
  _T_4726_im = _RAND_9059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9060 = {1{`RANDOM}};
  _T_4727_re = _RAND_9060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9061 = {1{`RANDOM}};
  _T_4727_im = _RAND_9061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9062 = {1{`RANDOM}};
  _T_4728_re = _RAND_9062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9063 = {1{`RANDOM}};
  _T_4728_im = _RAND_9063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9064 = {1{`RANDOM}};
  _T_4729_re = _RAND_9064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9065 = {1{`RANDOM}};
  _T_4729_im = _RAND_9065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9066 = {1{`RANDOM}};
  _T_4730_re = _RAND_9066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9067 = {1{`RANDOM}};
  _T_4730_im = _RAND_9067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9068 = {1{`RANDOM}};
  _T_4731_re = _RAND_9068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9069 = {1{`RANDOM}};
  _T_4731_im = _RAND_9069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9070 = {1{`RANDOM}};
  _T_4732_re = _RAND_9070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9071 = {1{`RANDOM}};
  _T_4732_im = _RAND_9071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9072 = {1{`RANDOM}};
  _T_4733_re = _RAND_9072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9073 = {1{`RANDOM}};
  _T_4733_im = _RAND_9073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9074 = {1{`RANDOM}};
  _T_4734_re = _RAND_9074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9075 = {1{`RANDOM}};
  _T_4734_im = _RAND_9075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9076 = {1{`RANDOM}};
  _T_4735_re = _RAND_9076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9077 = {1{`RANDOM}};
  _T_4735_im = _RAND_9077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9078 = {1{`RANDOM}};
  _T_4736_re = _RAND_9078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9079 = {1{`RANDOM}};
  _T_4736_im = _RAND_9079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9080 = {1{`RANDOM}};
  _T_4737_re = _RAND_9080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9081 = {1{`RANDOM}};
  _T_4737_im = _RAND_9081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9082 = {1{`RANDOM}};
  _T_4738_re = _RAND_9082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9083 = {1{`RANDOM}};
  _T_4738_im = _RAND_9083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9084 = {1{`RANDOM}};
  _T_4739_re = _RAND_9084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9085 = {1{`RANDOM}};
  _T_4739_im = _RAND_9085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9086 = {1{`RANDOM}};
  _T_4740_re = _RAND_9086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9087 = {1{`RANDOM}};
  _T_4740_im = _RAND_9087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9088 = {1{`RANDOM}};
  _T_4741_re = _RAND_9088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9089 = {1{`RANDOM}};
  _T_4741_im = _RAND_9089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9090 = {1{`RANDOM}};
  _T_4742_re = _RAND_9090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9091 = {1{`RANDOM}};
  _T_4742_im = _RAND_9091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9092 = {1{`RANDOM}};
  _T_4743_re = _RAND_9092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9093 = {1{`RANDOM}};
  _T_4743_im = _RAND_9093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9094 = {1{`RANDOM}};
  _T_4744_re = _RAND_9094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9095 = {1{`RANDOM}};
  _T_4744_im = _RAND_9095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9096 = {1{`RANDOM}};
  _T_4745_re = _RAND_9096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9097 = {1{`RANDOM}};
  _T_4745_im = _RAND_9097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9098 = {1{`RANDOM}};
  _T_4746_re = _RAND_9098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9099 = {1{`RANDOM}};
  _T_4746_im = _RAND_9099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9100 = {1{`RANDOM}};
  _T_4747_re = _RAND_9100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9101 = {1{`RANDOM}};
  _T_4747_im = _RAND_9101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9102 = {1{`RANDOM}};
  _T_4748_re = _RAND_9102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9103 = {1{`RANDOM}};
  _T_4748_im = _RAND_9103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9104 = {1{`RANDOM}};
  _T_4749_re = _RAND_9104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9105 = {1{`RANDOM}};
  _T_4749_im = _RAND_9105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9106 = {1{`RANDOM}};
  _T_4750_re = _RAND_9106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9107 = {1{`RANDOM}};
  _T_4750_im = _RAND_9107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9108 = {1{`RANDOM}};
  _T_4751_re = _RAND_9108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9109 = {1{`RANDOM}};
  _T_4751_im = _RAND_9109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9110 = {1{`RANDOM}};
  _T_4752_re = _RAND_9110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9111 = {1{`RANDOM}};
  _T_4752_im = _RAND_9111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9112 = {1{`RANDOM}};
  _T_4753_re = _RAND_9112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9113 = {1{`RANDOM}};
  _T_4753_im = _RAND_9113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9114 = {1{`RANDOM}};
  _T_4754_re = _RAND_9114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9115 = {1{`RANDOM}};
  _T_4754_im = _RAND_9115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9116 = {1{`RANDOM}};
  _T_4755_re = _RAND_9116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9117 = {1{`RANDOM}};
  _T_4755_im = _RAND_9117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9118 = {1{`RANDOM}};
  _T_4756_re = _RAND_9118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9119 = {1{`RANDOM}};
  _T_4756_im = _RAND_9119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9120 = {1{`RANDOM}};
  _T_4757_re = _RAND_9120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9121 = {1{`RANDOM}};
  _T_4757_im = _RAND_9121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9122 = {1{`RANDOM}};
  _T_4758_re = _RAND_9122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9123 = {1{`RANDOM}};
  _T_4758_im = _RAND_9123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9124 = {1{`RANDOM}};
  _T_4759_re = _RAND_9124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9125 = {1{`RANDOM}};
  _T_4759_im = _RAND_9125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9126 = {1{`RANDOM}};
  _T_4760_re = _RAND_9126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9127 = {1{`RANDOM}};
  _T_4760_im = _RAND_9127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9128 = {1{`RANDOM}};
  _T_4761_re = _RAND_9128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9129 = {1{`RANDOM}};
  _T_4761_im = _RAND_9129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9130 = {1{`RANDOM}};
  _T_4762_re = _RAND_9130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9131 = {1{`RANDOM}};
  _T_4762_im = _RAND_9131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9132 = {1{`RANDOM}};
  _T_4763_re = _RAND_9132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9133 = {1{`RANDOM}};
  _T_4763_im = _RAND_9133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9134 = {1{`RANDOM}};
  _T_4764_re = _RAND_9134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9135 = {1{`RANDOM}};
  _T_4764_im = _RAND_9135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9136 = {1{`RANDOM}};
  _T_4765_re = _RAND_9136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9137 = {1{`RANDOM}};
  _T_4765_im = _RAND_9137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9138 = {1{`RANDOM}};
  _T_4766_re = _RAND_9138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9139 = {1{`RANDOM}};
  _T_4766_im = _RAND_9139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9140 = {1{`RANDOM}};
  _T_4767_re = _RAND_9140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9141 = {1{`RANDOM}};
  _T_4767_im = _RAND_9141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9142 = {1{`RANDOM}};
  _T_4768_re = _RAND_9142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9143 = {1{`RANDOM}};
  _T_4768_im = _RAND_9143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9144 = {1{`RANDOM}};
  _T_4769_re = _RAND_9144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9145 = {1{`RANDOM}};
  _T_4769_im = _RAND_9145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9146 = {1{`RANDOM}};
  _T_4770_re = _RAND_9146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9147 = {1{`RANDOM}};
  _T_4770_im = _RAND_9147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9148 = {1{`RANDOM}};
  _T_4771_re = _RAND_9148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9149 = {1{`RANDOM}};
  _T_4771_im = _RAND_9149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9150 = {1{`RANDOM}};
  _T_4772_re = _RAND_9150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9151 = {1{`RANDOM}};
  _T_4772_im = _RAND_9151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9152 = {1{`RANDOM}};
  _T_4773_re = _RAND_9152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9153 = {1{`RANDOM}};
  _T_4773_im = _RAND_9153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9154 = {1{`RANDOM}};
  _T_4774_re = _RAND_9154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9155 = {1{`RANDOM}};
  _T_4774_im = _RAND_9155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9156 = {1{`RANDOM}};
  _T_4775_re = _RAND_9156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9157 = {1{`RANDOM}};
  _T_4775_im = _RAND_9157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9158 = {1{`RANDOM}};
  _T_4776_re = _RAND_9158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9159 = {1{`RANDOM}};
  _T_4776_im = _RAND_9159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9160 = {1{`RANDOM}};
  _T_4777_re = _RAND_9160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9161 = {1{`RANDOM}};
  _T_4777_im = _RAND_9161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9162 = {1{`RANDOM}};
  _T_4778_re = _RAND_9162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9163 = {1{`RANDOM}};
  _T_4778_im = _RAND_9163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9164 = {1{`RANDOM}};
  _T_4779_re = _RAND_9164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9165 = {1{`RANDOM}};
  _T_4779_im = _RAND_9165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9166 = {1{`RANDOM}};
  _T_4780_re = _RAND_9166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9167 = {1{`RANDOM}};
  _T_4780_im = _RAND_9167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9168 = {1{`RANDOM}};
  _T_4781_re = _RAND_9168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9169 = {1{`RANDOM}};
  _T_4781_im = _RAND_9169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9170 = {1{`RANDOM}};
  _T_4782_re = _RAND_9170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9171 = {1{`RANDOM}};
  _T_4782_im = _RAND_9171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9172 = {1{`RANDOM}};
  _T_4783_re = _RAND_9172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9173 = {1{`RANDOM}};
  _T_4783_im = _RAND_9173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9174 = {1{`RANDOM}};
  _T_4784_re = _RAND_9174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9175 = {1{`RANDOM}};
  _T_4784_im = _RAND_9175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9176 = {1{`RANDOM}};
  _T_4785_re = _RAND_9176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9177 = {1{`RANDOM}};
  _T_4785_im = _RAND_9177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9178 = {1{`RANDOM}};
  _T_4786_re = _RAND_9178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9179 = {1{`RANDOM}};
  _T_4786_im = _RAND_9179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9180 = {1{`RANDOM}};
  _T_4787_re = _RAND_9180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9181 = {1{`RANDOM}};
  _T_4787_im = _RAND_9181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9182 = {1{`RANDOM}};
  _T_4788_re = _RAND_9182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9183 = {1{`RANDOM}};
  _T_4788_im = _RAND_9183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9184 = {1{`RANDOM}};
  _T_4789_re = _RAND_9184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9185 = {1{`RANDOM}};
  _T_4789_im = _RAND_9185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9186 = {1{`RANDOM}};
  _T_4790_re = _RAND_9186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9187 = {1{`RANDOM}};
  _T_4790_im = _RAND_9187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9188 = {1{`RANDOM}};
  _T_4791_re = _RAND_9188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9189 = {1{`RANDOM}};
  _T_4791_im = _RAND_9189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9190 = {1{`RANDOM}};
  _T_4792_re = _RAND_9190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9191 = {1{`RANDOM}};
  _T_4792_im = _RAND_9191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9192 = {1{`RANDOM}};
  _T_4793_re = _RAND_9192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9193 = {1{`RANDOM}};
  _T_4793_im = _RAND_9193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9194 = {1{`RANDOM}};
  _T_4794_re = _RAND_9194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9195 = {1{`RANDOM}};
  _T_4794_im = _RAND_9195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9196 = {1{`RANDOM}};
  _T_4795_re = _RAND_9196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9197 = {1{`RANDOM}};
  _T_4795_im = _RAND_9197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9198 = {1{`RANDOM}};
  _T_4796_re = _RAND_9198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9199 = {1{`RANDOM}};
  _T_4796_im = _RAND_9199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9200 = {1{`RANDOM}};
  _T_4797_re = _RAND_9200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9201 = {1{`RANDOM}};
  _T_4797_im = _RAND_9201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9202 = {1{`RANDOM}};
  _T_4798_re = _RAND_9202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9203 = {1{`RANDOM}};
  _T_4798_im = _RAND_9203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9204 = {1{`RANDOM}};
  _T_4799_re = _RAND_9204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9205 = {1{`RANDOM}};
  _T_4799_im = _RAND_9205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9206 = {1{`RANDOM}};
  _T_4800_re = _RAND_9206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9207 = {1{`RANDOM}};
  _T_4800_im = _RAND_9207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9208 = {1{`RANDOM}};
  _T_4801_re = _RAND_9208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9209 = {1{`RANDOM}};
  _T_4801_im = _RAND_9209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9210 = {1{`RANDOM}};
  _T_4802_re = _RAND_9210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9211 = {1{`RANDOM}};
  _T_4802_im = _RAND_9211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9212 = {1{`RANDOM}};
  _T_4803_re = _RAND_9212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9213 = {1{`RANDOM}};
  _T_4803_im = _RAND_9213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9214 = {1{`RANDOM}};
  _T_4804_re = _RAND_9214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9215 = {1{`RANDOM}};
  _T_4804_im = _RAND_9215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9216 = {1{`RANDOM}};
  _T_4805_re = _RAND_9216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9217 = {1{`RANDOM}};
  _T_4805_im = _RAND_9217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9218 = {1{`RANDOM}};
  _T_4811_re = _RAND_9218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9219 = {1{`RANDOM}};
  _T_4811_im = _RAND_9219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9220 = {1{`RANDOM}};
  _T_4812_re = _RAND_9220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9221 = {1{`RANDOM}};
  _T_4812_im = _RAND_9221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9222 = {1{`RANDOM}};
  _T_4813_re = _RAND_9222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9223 = {1{`RANDOM}};
  _T_4813_im = _RAND_9223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9224 = {1{`RANDOM}};
  _T_4814_re = _RAND_9224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9225 = {1{`RANDOM}};
  _T_4814_im = _RAND_9225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9226 = {1{`RANDOM}};
  _T_4815_re = _RAND_9226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9227 = {1{`RANDOM}};
  _T_4815_im = _RAND_9227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9228 = {1{`RANDOM}};
  _T_4816_re = _RAND_9228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9229 = {1{`RANDOM}};
  _T_4816_im = _RAND_9229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9230 = {1{`RANDOM}};
  _T_4817_re = _RAND_9230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9231 = {1{`RANDOM}};
  _T_4817_im = _RAND_9231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9232 = {1{`RANDOM}};
  _T_4818_re = _RAND_9232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9233 = {1{`RANDOM}};
  _T_4818_im = _RAND_9233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9234 = {1{`RANDOM}};
  _T_4819_re = _RAND_9234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9235 = {1{`RANDOM}};
  _T_4819_im = _RAND_9235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9236 = {1{`RANDOM}};
  _T_4820_re = _RAND_9236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9237 = {1{`RANDOM}};
  _T_4820_im = _RAND_9237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9238 = {1{`RANDOM}};
  _T_4821_re = _RAND_9238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9239 = {1{`RANDOM}};
  _T_4821_im = _RAND_9239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9240 = {1{`RANDOM}};
  _T_4822_re = _RAND_9240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9241 = {1{`RANDOM}};
  _T_4822_im = _RAND_9241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9242 = {1{`RANDOM}};
  _T_4823_re = _RAND_9242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9243 = {1{`RANDOM}};
  _T_4823_im = _RAND_9243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9244 = {1{`RANDOM}};
  _T_4824_re = _RAND_9244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9245 = {1{`RANDOM}};
  _T_4824_im = _RAND_9245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9246 = {1{`RANDOM}};
  _T_4825_re = _RAND_9246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9247 = {1{`RANDOM}};
  _T_4825_im = _RAND_9247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9248 = {1{`RANDOM}};
  _T_4826_re = _RAND_9248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9249 = {1{`RANDOM}};
  _T_4826_im = _RAND_9249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9250 = {1{`RANDOM}};
  _T_4827_re = _RAND_9250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9251 = {1{`RANDOM}};
  _T_4827_im = _RAND_9251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9252 = {1{`RANDOM}};
  _T_4828_re = _RAND_9252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9253 = {1{`RANDOM}};
  _T_4828_im = _RAND_9253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9254 = {1{`RANDOM}};
  _T_4829_re = _RAND_9254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9255 = {1{`RANDOM}};
  _T_4829_im = _RAND_9255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9256 = {1{`RANDOM}};
  _T_4830_re = _RAND_9256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9257 = {1{`RANDOM}};
  _T_4830_im = _RAND_9257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9258 = {1{`RANDOM}};
  _T_4831_re = _RAND_9258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9259 = {1{`RANDOM}};
  _T_4831_im = _RAND_9259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9260 = {1{`RANDOM}};
  _T_4832_re = _RAND_9260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9261 = {1{`RANDOM}};
  _T_4832_im = _RAND_9261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9262 = {1{`RANDOM}};
  _T_4833_re = _RAND_9262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9263 = {1{`RANDOM}};
  _T_4833_im = _RAND_9263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9264 = {1{`RANDOM}};
  _T_4834_re = _RAND_9264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9265 = {1{`RANDOM}};
  _T_4834_im = _RAND_9265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9266 = {1{`RANDOM}};
  _T_4835_re = _RAND_9266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9267 = {1{`RANDOM}};
  _T_4835_im = _RAND_9267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9268 = {1{`RANDOM}};
  _T_4836_re = _RAND_9268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9269 = {1{`RANDOM}};
  _T_4836_im = _RAND_9269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9270 = {1{`RANDOM}};
  _T_4837_re = _RAND_9270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9271 = {1{`RANDOM}};
  _T_4837_im = _RAND_9271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9272 = {1{`RANDOM}};
  _T_4838_re = _RAND_9272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9273 = {1{`RANDOM}};
  _T_4838_im = _RAND_9273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9274 = {1{`RANDOM}};
  _T_4839_re = _RAND_9274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9275 = {1{`RANDOM}};
  _T_4839_im = _RAND_9275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9276 = {1{`RANDOM}};
  _T_4840_re = _RAND_9276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9277 = {1{`RANDOM}};
  _T_4840_im = _RAND_9277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9278 = {1{`RANDOM}};
  _T_4841_re = _RAND_9278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9279 = {1{`RANDOM}};
  _T_4841_im = _RAND_9279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9280 = {1{`RANDOM}};
  _T_4842_re = _RAND_9280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9281 = {1{`RANDOM}};
  _T_4842_im = _RAND_9281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9282 = {1{`RANDOM}};
  _T_4843_re = _RAND_9282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9283 = {1{`RANDOM}};
  _T_4843_im = _RAND_9283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9284 = {1{`RANDOM}};
  _T_4844_re = _RAND_9284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9285 = {1{`RANDOM}};
  _T_4844_im = _RAND_9285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9286 = {1{`RANDOM}};
  _T_4845_re = _RAND_9286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9287 = {1{`RANDOM}};
  _T_4845_im = _RAND_9287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9288 = {1{`RANDOM}};
  _T_4846_re = _RAND_9288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9289 = {1{`RANDOM}};
  _T_4846_im = _RAND_9289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9290 = {1{`RANDOM}};
  _T_4847_re = _RAND_9290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9291 = {1{`RANDOM}};
  _T_4847_im = _RAND_9291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9292 = {1{`RANDOM}};
  _T_4848_re = _RAND_9292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9293 = {1{`RANDOM}};
  _T_4848_im = _RAND_9293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9294 = {1{`RANDOM}};
  _T_4849_re = _RAND_9294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9295 = {1{`RANDOM}};
  _T_4849_im = _RAND_9295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9296 = {1{`RANDOM}};
  _T_4850_re = _RAND_9296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9297 = {1{`RANDOM}};
  _T_4850_im = _RAND_9297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9298 = {1{`RANDOM}};
  _T_4851_re = _RAND_9298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9299 = {1{`RANDOM}};
  _T_4851_im = _RAND_9299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9300 = {1{`RANDOM}};
  _T_4852_re = _RAND_9300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9301 = {1{`RANDOM}};
  _T_4852_im = _RAND_9301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9302 = {1{`RANDOM}};
  _T_4853_re = _RAND_9302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9303 = {1{`RANDOM}};
  _T_4853_im = _RAND_9303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9304 = {1{`RANDOM}};
  _T_4854_re = _RAND_9304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9305 = {1{`RANDOM}};
  _T_4854_im = _RAND_9305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9306 = {1{`RANDOM}};
  _T_4855_re = _RAND_9306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9307 = {1{`RANDOM}};
  _T_4855_im = _RAND_9307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9308 = {1{`RANDOM}};
  _T_4856_re = _RAND_9308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9309 = {1{`RANDOM}};
  _T_4856_im = _RAND_9309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9310 = {1{`RANDOM}};
  _T_4857_re = _RAND_9310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9311 = {1{`RANDOM}};
  _T_4857_im = _RAND_9311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9312 = {1{`RANDOM}};
  _T_4858_re = _RAND_9312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9313 = {1{`RANDOM}};
  _T_4858_im = _RAND_9313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9314 = {1{`RANDOM}};
  _T_4859_re = _RAND_9314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9315 = {1{`RANDOM}};
  _T_4859_im = _RAND_9315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9316 = {1{`RANDOM}};
  _T_4860_re = _RAND_9316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9317 = {1{`RANDOM}};
  _T_4860_im = _RAND_9317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9318 = {1{`RANDOM}};
  _T_4861_re = _RAND_9318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9319 = {1{`RANDOM}};
  _T_4861_im = _RAND_9319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9320 = {1{`RANDOM}};
  _T_4862_re = _RAND_9320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9321 = {1{`RANDOM}};
  _T_4862_im = _RAND_9321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9322 = {1{`RANDOM}};
  _T_4863_re = _RAND_9322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9323 = {1{`RANDOM}};
  _T_4863_im = _RAND_9323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9324 = {1{`RANDOM}};
  _T_4864_re = _RAND_9324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9325 = {1{`RANDOM}};
  _T_4864_im = _RAND_9325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9326 = {1{`RANDOM}};
  _T_4865_re = _RAND_9326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9327 = {1{`RANDOM}};
  _T_4865_im = _RAND_9327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9328 = {1{`RANDOM}};
  _T_4866_re = _RAND_9328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9329 = {1{`RANDOM}};
  _T_4866_im = _RAND_9329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9330 = {1{`RANDOM}};
  _T_4867_re = _RAND_9330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9331 = {1{`RANDOM}};
  _T_4867_im = _RAND_9331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9332 = {1{`RANDOM}};
  _T_4868_re = _RAND_9332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9333 = {1{`RANDOM}};
  _T_4868_im = _RAND_9333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9334 = {1{`RANDOM}};
  _T_4869_re = _RAND_9334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9335 = {1{`RANDOM}};
  _T_4869_im = _RAND_9335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9336 = {1{`RANDOM}};
  _T_4870_re = _RAND_9336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9337 = {1{`RANDOM}};
  _T_4870_im = _RAND_9337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9338 = {1{`RANDOM}};
  _T_4871_re = _RAND_9338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9339 = {1{`RANDOM}};
  _T_4871_im = _RAND_9339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9340 = {1{`RANDOM}};
  _T_4872_re = _RAND_9340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9341 = {1{`RANDOM}};
  _T_4872_im = _RAND_9341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9342 = {1{`RANDOM}};
  _T_4873_re = _RAND_9342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9343 = {1{`RANDOM}};
  _T_4873_im = _RAND_9343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9344 = {1{`RANDOM}};
  _T_4874_re = _RAND_9344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9345 = {1{`RANDOM}};
  _T_4874_im = _RAND_9345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9346 = {1{`RANDOM}};
  _T_4875_re = _RAND_9346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9347 = {1{`RANDOM}};
  _T_4875_im = _RAND_9347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9348 = {1{`RANDOM}};
  _T_4876_re = _RAND_9348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9349 = {1{`RANDOM}};
  _T_4876_im = _RAND_9349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9350 = {1{`RANDOM}};
  _T_4877_re = _RAND_9350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9351 = {1{`RANDOM}};
  _T_4877_im = _RAND_9351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9352 = {1{`RANDOM}};
  _T_4878_re = _RAND_9352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9353 = {1{`RANDOM}};
  _T_4878_im = _RAND_9353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9354 = {1{`RANDOM}};
  _T_4879_re = _RAND_9354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9355 = {1{`RANDOM}};
  _T_4879_im = _RAND_9355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9356 = {1{`RANDOM}};
  _T_4880_re = _RAND_9356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9357 = {1{`RANDOM}};
  _T_4880_im = _RAND_9357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9358 = {1{`RANDOM}};
  _T_4881_re = _RAND_9358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9359 = {1{`RANDOM}};
  _T_4881_im = _RAND_9359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9360 = {1{`RANDOM}};
  _T_4882_re = _RAND_9360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9361 = {1{`RANDOM}};
  _T_4882_im = _RAND_9361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9362 = {1{`RANDOM}};
  _T_4883_re = _RAND_9362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9363 = {1{`RANDOM}};
  _T_4883_im = _RAND_9363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9364 = {1{`RANDOM}};
  _T_4884_re = _RAND_9364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9365 = {1{`RANDOM}};
  _T_4884_im = _RAND_9365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9366 = {1{`RANDOM}};
  _T_4885_re = _RAND_9366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9367 = {1{`RANDOM}};
  _T_4885_im = _RAND_9367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9368 = {1{`RANDOM}};
  _T_4886_re = _RAND_9368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9369 = {1{`RANDOM}};
  _T_4886_im = _RAND_9369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9370 = {1{`RANDOM}};
  _T_4887_re = _RAND_9370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9371 = {1{`RANDOM}};
  _T_4887_im = _RAND_9371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9372 = {1{`RANDOM}};
  _T_4888_re = _RAND_9372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9373 = {1{`RANDOM}};
  _T_4888_im = _RAND_9373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9374 = {1{`RANDOM}};
  _T_4889_re = _RAND_9374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9375 = {1{`RANDOM}};
  _T_4889_im = _RAND_9375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9376 = {1{`RANDOM}};
  _T_4890_re = _RAND_9376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9377 = {1{`RANDOM}};
  _T_4890_im = _RAND_9377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9378 = {1{`RANDOM}};
  _T_4891_re = _RAND_9378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9379 = {1{`RANDOM}};
  _T_4891_im = _RAND_9379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9380 = {1{`RANDOM}};
  _T_4892_re = _RAND_9380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9381 = {1{`RANDOM}};
  _T_4892_im = _RAND_9381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9382 = {1{`RANDOM}};
  _T_4893_re = _RAND_9382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9383 = {1{`RANDOM}};
  _T_4893_im = _RAND_9383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9384 = {1{`RANDOM}};
  _T_4894_re = _RAND_9384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9385 = {1{`RANDOM}};
  _T_4894_im = _RAND_9385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9386 = {1{`RANDOM}};
  _T_4895_re = _RAND_9386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9387 = {1{`RANDOM}};
  _T_4895_im = _RAND_9387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9388 = {1{`RANDOM}};
  _T_4896_re = _RAND_9388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9389 = {1{`RANDOM}};
  _T_4896_im = _RAND_9389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9390 = {1{`RANDOM}};
  _T_4897_re = _RAND_9390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9391 = {1{`RANDOM}};
  _T_4897_im = _RAND_9391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9392 = {1{`RANDOM}};
  _T_4898_re = _RAND_9392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9393 = {1{`RANDOM}};
  _T_4898_im = _RAND_9393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9394 = {1{`RANDOM}};
  _T_4899_re = _RAND_9394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9395 = {1{`RANDOM}};
  _T_4899_im = _RAND_9395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9396 = {1{`RANDOM}};
  _T_4900_re = _RAND_9396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9397 = {1{`RANDOM}};
  _T_4900_im = _RAND_9397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9398 = {1{`RANDOM}};
  _T_4901_re = _RAND_9398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9399 = {1{`RANDOM}};
  _T_4901_im = _RAND_9399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9400 = {1{`RANDOM}};
  _T_4902_re = _RAND_9400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9401 = {1{`RANDOM}};
  _T_4902_im = _RAND_9401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9402 = {1{`RANDOM}};
  _T_4903_re = _RAND_9402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9403 = {1{`RANDOM}};
  _T_4903_im = _RAND_9403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9404 = {1{`RANDOM}};
  _T_4904_re = _RAND_9404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9405 = {1{`RANDOM}};
  _T_4904_im = _RAND_9405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9406 = {1{`RANDOM}};
  _T_4905_re = _RAND_9406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9407 = {1{`RANDOM}};
  _T_4905_im = _RAND_9407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9408 = {1{`RANDOM}};
  _T_4906_re = _RAND_9408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9409 = {1{`RANDOM}};
  _T_4906_im = _RAND_9409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9410 = {1{`RANDOM}};
  _T_4907_re = _RAND_9410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9411 = {1{`RANDOM}};
  _T_4907_im = _RAND_9411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9412 = {1{`RANDOM}};
  _T_4908_re = _RAND_9412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9413 = {1{`RANDOM}};
  _T_4908_im = _RAND_9413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9414 = {1{`RANDOM}};
  _T_4909_re = _RAND_9414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9415 = {1{`RANDOM}};
  _T_4909_im = _RAND_9415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9416 = {1{`RANDOM}};
  _T_4910_re = _RAND_9416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9417 = {1{`RANDOM}};
  _T_4910_im = _RAND_9417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9418 = {1{`RANDOM}};
  _T_4911_re = _RAND_9418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9419 = {1{`RANDOM}};
  _T_4911_im = _RAND_9419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9420 = {1{`RANDOM}};
  _T_4912_re = _RAND_9420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9421 = {1{`RANDOM}};
  _T_4912_im = _RAND_9421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9422 = {1{`RANDOM}};
  _T_4913_re = _RAND_9422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9423 = {1{`RANDOM}};
  _T_4913_im = _RAND_9423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9424 = {1{`RANDOM}};
  _T_4914_re = _RAND_9424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9425 = {1{`RANDOM}};
  _T_4914_im = _RAND_9425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9426 = {1{`RANDOM}};
  _T_4915_re = _RAND_9426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9427 = {1{`RANDOM}};
  _T_4915_im = _RAND_9427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9428 = {1{`RANDOM}};
  _T_4916_re = _RAND_9428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9429 = {1{`RANDOM}};
  _T_4916_im = _RAND_9429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9430 = {1{`RANDOM}};
  _T_4917_re = _RAND_9430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9431 = {1{`RANDOM}};
  _T_4917_im = _RAND_9431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9432 = {1{`RANDOM}};
  _T_4918_re = _RAND_9432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9433 = {1{`RANDOM}};
  _T_4918_im = _RAND_9433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9434 = {1{`RANDOM}};
  _T_4919_re = _RAND_9434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9435 = {1{`RANDOM}};
  _T_4919_im = _RAND_9435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9436 = {1{`RANDOM}};
  _T_4920_re = _RAND_9436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9437 = {1{`RANDOM}};
  _T_4920_im = _RAND_9437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9438 = {1{`RANDOM}};
  _T_4921_re = _RAND_9438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9439 = {1{`RANDOM}};
  _T_4921_im = _RAND_9439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9440 = {1{`RANDOM}};
  _T_4922_re = _RAND_9440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9441 = {1{`RANDOM}};
  _T_4922_im = _RAND_9441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9442 = {1{`RANDOM}};
  _T_4923_re = _RAND_9442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9443 = {1{`RANDOM}};
  _T_4923_im = _RAND_9443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9444 = {1{`RANDOM}};
  _T_4924_re = _RAND_9444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9445 = {1{`RANDOM}};
  _T_4924_im = _RAND_9445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9446 = {1{`RANDOM}};
  _T_4925_re = _RAND_9446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9447 = {1{`RANDOM}};
  _T_4925_im = _RAND_9447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9448 = {1{`RANDOM}};
  _T_4926_re = _RAND_9448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9449 = {1{`RANDOM}};
  _T_4926_im = _RAND_9449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9450 = {1{`RANDOM}};
  _T_4927_re = _RAND_9450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9451 = {1{`RANDOM}};
  _T_4927_im = _RAND_9451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9452 = {1{`RANDOM}};
  _T_4928_re = _RAND_9452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9453 = {1{`RANDOM}};
  _T_4928_im = _RAND_9453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9454 = {1{`RANDOM}};
  _T_4929_re = _RAND_9454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9455 = {1{`RANDOM}};
  _T_4929_im = _RAND_9455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9456 = {1{`RANDOM}};
  _T_4930_re = _RAND_9456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9457 = {1{`RANDOM}};
  _T_4930_im = _RAND_9457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9458 = {1{`RANDOM}};
  _T_4931_re = _RAND_9458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9459 = {1{`RANDOM}};
  _T_4931_im = _RAND_9459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9460 = {1{`RANDOM}};
  _T_4932_re = _RAND_9460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9461 = {1{`RANDOM}};
  _T_4932_im = _RAND_9461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9462 = {1{`RANDOM}};
  _T_4933_re = _RAND_9462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9463 = {1{`RANDOM}};
  _T_4933_im = _RAND_9463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9464 = {1{`RANDOM}};
  _T_4934_re = _RAND_9464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9465 = {1{`RANDOM}};
  _T_4934_im = _RAND_9465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9466 = {1{`RANDOM}};
  _T_4935_re = _RAND_9466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9467 = {1{`RANDOM}};
  _T_4935_im = _RAND_9467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9468 = {1{`RANDOM}};
  _T_4936_re = _RAND_9468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9469 = {1{`RANDOM}};
  _T_4936_im = _RAND_9469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9470 = {1{`RANDOM}};
  _T_4937_re = _RAND_9470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9471 = {1{`RANDOM}};
  _T_4937_im = _RAND_9471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9472 = {1{`RANDOM}};
  _T_4938_re = _RAND_9472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9473 = {1{`RANDOM}};
  _T_4938_im = _RAND_9473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9474 = {1{`RANDOM}};
  _T_4939_re = _RAND_9474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9475 = {1{`RANDOM}};
  _T_4939_im = _RAND_9475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9476 = {1{`RANDOM}};
  _T_4940_re = _RAND_9476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9477 = {1{`RANDOM}};
  _T_4940_im = _RAND_9477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9478 = {1{`RANDOM}};
  _T_4941_re = _RAND_9478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9479 = {1{`RANDOM}};
  _T_4941_im = _RAND_9479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9480 = {1{`RANDOM}};
  _T_4942_re = _RAND_9480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9481 = {1{`RANDOM}};
  _T_4942_im = _RAND_9481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9482 = {1{`RANDOM}};
  _T_4943_re = _RAND_9482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9483 = {1{`RANDOM}};
  _T_4943_im = _RAND_9483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9484 = {1{`RANDOM}};
  _T_4944_re = _RAND_9484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9485 = {1{`RANDOM}};
  _T_4944_im = _RAND_9485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9486 = {1{`RANDOM}};
  _T_4945_re = _RAND_9486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9487 = {1{`RANDOM}};
  _T_4945_im = _RAND_9487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9488 = {1{`RANDOM}};
  _T_4946_re = _RAND_9488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9489 = {1{`RANDOM}};
  _T_4946_im = _RAND_9489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9490 = {1{`RANDOM}};
  _T_4947_re = _RAND_9490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9491 = {1{`RANDOM}};
  _T_4947_im = _RAND_9491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9492 = {1{`RANDOM}};
  _T_4948_re = _RAND_9492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9493 = {1{`RANDOM}};
  _T_4948_im = _RAND_9493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9494 = {1{`RANDOM}};
  _T_4949_re = _RAND_9494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9495 = {1{`RANDOM}};
  _T_4949_im = _RAND_9495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9496 = {1{`RANDOM}};
  _T_4950_re = _RAND_9496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9497 = {1{`RANDOM}};
  _T_4950_im = _RAND_9497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9498 = {1{`RANDOM}};
  _T_4951_re = _RAND_9498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9499 = {1{`RANDOM}};
  _T_4951_im = _RAND_9499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9500 = {1{`RANDOM}};
  _T_4952_re = _RAND_9500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9501 = {1{`RANDOM}};
  _T_4952_im = _RAND_9501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9502 = {1{`RANDOM}};
  _T_4953_re = _RAND_9502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9503 = {1{`RANDOM}};
  _T_4953_im = _RAND_9503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9504 = {1{`RANDOM}};
  _T_4954_re = _RAND_9504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9505 = {1{`RANDOM}};
  _T_4954_im = _RAND_9505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9506 = {1{`RANDOM}};
  _T_4955_re = _RAND_9506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9507 = {1{`RANDOM}};
  _T_4955_im = _RAND_9507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9508 = {1{`RANDOM}};
  _T_4956_re = _RAND_9508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9509 = {1{`RANDOM}};
  _T_4956_im = _RAND_9509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9510 = {1{`RANDOM}};
  _T_4957_re = _RAND_9510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9511 = {1{`RANDOM}};
  _T_4957_im = _RAND_9511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9512 = {1{`RANDOM}};
  _T_4958_re = _RAND_9512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9513 = {1{`RANDOM}};
  _T_4958_im = _RAND_9513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9514 = {1{`RANDOM}};
  _T_4959_re = _RAND_9514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9515 = {1{`RANDOM}};
  _T_4959_im = _RAND_9515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9516 = {1{`RANDOM}};
  _T_4960_re = _RAND_9516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9517 = {1{`RANDOM}};
  _T_4960_im = _RAND_9517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9518 = {1{`RANDOM}};
  _T_4961_re = _RAND_9518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9519 = {1{`RANDOM}};
  _T_4961_im = _RAND_9519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9520 = {1{`RANDOM}};
  _T_4962_re = _RAND_9520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9521 = {1{`RANDOM}};
  _T_4962_im = _RAND_9521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9522 = {1{`RANDOM}};
  _T_4963_re = _RAND_9522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9523 = {1{`RANDOM}};
  _T_4963_im = _RAND_9523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9524 = {1{`RANDOM}};
  _T_4964_re = _RAND_9524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9525 = {1{`RANDOM}};
  _T_4964_im = _RAND_9525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9526 = {1{`RANDOM}};
  _T_4965_re = _RAND_9526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9527 = {1{`RANDOM}};
  _T_4965_im = _RAND_9527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9528 = {1{`RANDOM}};
  _T_4966_re = _RAND_9528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9529 = {1{`RANDOM}};
  _T_4966_im = _RAND_9529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9530 = {1{`RANDOM}};
  _T_4967_re = _RAND_9530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9531 = {1{`RANDOM}};
  _T_4967_im = _RAND_9531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9532 = {1{`RANDOM}};
  _T_4968_re = _RAND_9532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9533 = {1{`RANDOM}};
  _T_4968_im = _RAND_9533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9534 = {1{`RANDOM}};
  _T_4969_re = _RAND_9534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9535 = {1{`RANDOM}};
  _T_4969_im = _RAND_9535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9536 = {1{`RANDOM}};
  _T_4970_re = _RAND_9536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9537 = {1{`RANDOM}};
  _T_4970_im = _RAND_9537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9538 = {1{`RANDOM}};
  _T_4971_re = _RAND_9538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9539 = {1{`RANDOM}};
  _T_4971_im = _RAND_9539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9540 = {1{`RANDOM}};
  _T_4972_re = _RAND_9540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9541 = {1{`RANDOM}};
  _T_4972_im = _RAND_9541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9542 = {1{`RANDOM}};
  _T_4973_re = _RAND_9542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9543 = {1{`RANDOM}};
  _T_4973_im = _RAND_9543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9544 = {1{`RANDOM}};
  _T_4974_re = _RAND_9544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9545 = {1{`RANDOM}};
  _T_4974_im = _RAND_9545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9546 = {1{`RANDOM}};
  _T_4975_re = _RAND_9546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9547 = {1{`RANDOM}};
  _T_4975_im = _RAND_9547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9548 = {1{`RANDOM}};
  _T_4976_re = _RAND_9548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9549 = {1{`RANDOM}};
  _T_4976_im = _RAND_9549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9550 = {1{`RANDOM}};
  _T_4977_re = _RAND_9550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9551 = {1{`RANDOM}};
  _T_4977_im = _RAND_9551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9552 = {1{`RANDOM}};
  _T_4978_re = _RAND_9552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9553 = {1{`RANDOM}};
  _T_4978_im = _RAND_9553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9554 = {1{`RANDOM}};
  _T_4979_re = _RAND_9554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9555 = {1{`RANDOM}};
  _T_4979_im = _RAND_9555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9556 = {1{`RANDOM}};
  _T_4980_re = _RAND_9556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9557 = {1{`RANDOM}};
  _T_4980_im = _RAND_9557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9558 = {1{`RANDOM}};
  _T_4981_re = _RAND_9558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9559 = {1{`RANDOM}};
  _T_4981_im = _RAND_9559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9560 = {1{`RANDOM}};
  _T_4982_re = _RAND_9560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9561 = {1{`RANDOM}};
  _T_4982_im = _RAND_9561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9562 = {1{`RANDOM}};
  _T_4983_re = _RAND_9562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9563 = {1{`RANDOM}};
  _T_4983_im = _RAND_9563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9564 = {1{`RANDOM}};
  _T_4984_re = _RAND_9564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9565 = {1{`RANDOM}};
  _T_4984_im = _RAND_9565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9566 = {1{`RANDOM}};
  _T_4985_re = _RAND_9566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9567 = {1{`RANDOM}};
  _T_4985_im = _RAND_9567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9568 = {1{`RANDOM}};
  _T_4986_re = _RAND_9568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9569 = {1{`RANDOM}};
  _T_4986_im = _RAND_9569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9570 = {1{`RANDOM}};
  _T_4987_re = _RAND_9570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9571 = {1{`RANDOM}};
  _T_4987_im = _RAND_9571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9572 = {1{`RANDOM}};
  _T_4988_re = _RAND_9572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9573 = {1{`RANDOM}};
  _T_4988_im = _RAND_9573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9574 = {1{`RANDOM}};
  _T_4989_re = _RAND_9574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9575 = {1{`RANDOM}};
  _T_4989_im = _RAND_9575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9576 = {1{`RANDOM}};
  _T_4990_re = _RAND_9576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9577 = {1{`RANDOM}};
  _T_4990_im = _RAND_9577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9578 = {1{`RANDOM}};
  _T_4991_re = _RAND_9578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9579 = {1{`RANDOM}};
  _T_4991_im = _RAND_9579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9580 = {1{`RANDOM}};
  _T_4992_re = _RAND_9580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9581 = {1{`RANDOM}};
  _T_4992_im = _RAND_9581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9582 = {1{`RANDOM}};
  _T_4993_re = _RAND_9582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9583 = {1{`RANDOM}};
  _T_4993_im = _RAND_9583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9584 = {1{`RANDOM}};
  _T_4994_re = _RAND_9584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9585 = {1{`RANDOM}};
  _T_4994_im = _RAND_9585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9586 = {1{`RANDOM}};
  _T_4995_re = _RAND_9586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9587 = {1{`RANDOM}};
  _T_4995_im = _RAND_9587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9588 = {1{`RANDOM}};
  _T_4996_re = _RAND_9588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9589 = {1{`RANDOM}};
  _T_4996_im = _RAND_9589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9590 = {1{`RANDOM}};
  _T_4997_re = _RAND_9590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9591 = {1{`RANDOM}};
  _T_4997_im = _RAND_9591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9592 = {1{`RANDOM}};
  _T_4998_re = _RAND_9592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9593 = {1{`RANDOM}};
  _T_4998_im = _RAND_9593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9594 = {1{`RANDOM}};
  _T_4999_re = _RAND_9594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9595 = {1{`RANDOM}};
  _T_4999_im = _RAND_9595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9596 = {1{`RANDOM}};
  _T_5000_re = _RAND_9596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9597 = {1{`RANDOM}};
  _T_5000_im = _RAND_9597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9598 = {1{`RANDOM}};
  _T_5001_re = _RAND_9598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9599 = {1{`RANDOM}};
  _T_5001_im = _RAND_9599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9600 = {1{`RANDOM}};
  _T_5002_re = _RAND_9600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9601 = {1{`RANDOM}};
  _T_5002_im = _RAND_9601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9602 = {1{`RANDOM}};
  _T_5003_re = _RAND_9602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9603 = {1{`RANDOM}};
  _T_5003_im = _RAND_9603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9604 = {1{`RANDOM}};
  _T_5004_re = _RAND_9604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9605 = {1{`RANDOM}};
  _T_5004_im = _RAND_9605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9606 = {1{`RANDOM}};
  _T_5005_re = _RAND_9606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9607 = {1{`RANDOM}};
  _T_5005_im = _RAND_9607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9608 = {1{`RANDOM}};
  _T_5006_re = _RAND_9608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9609 = {1{`RANDOM}};
  _T_5006_im = _RAND_9609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9610 = {1{`RANDOM}};
  _T_5007_re = _RAND_9610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9611 = {1{`RANDOM}};
  _T_5007_im = _RAND_9611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9612 = {1{`RANDOM}};
  _T_5008_re = _RAND_9612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9613 = {1{`RANDOM}};
  _T_5008_im = _RAND_9613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9614 = {1{`RANDOM}};
  _T_5009_re = _RAND_9614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9615 = {1{`RANDOM}};
  _T_5009_im = _RAND_9615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9616 = {1{`RANDOM}};
  _T_5010_re = _RAND_9616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9617 = {1{`RANDOM}};
  _T_5010_im = _RAND_9617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9618 = {1{`RANDOM}};
  _T_5011_re = _RAND_9618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9619 = {1{`RANDOM}};
  _T_5011_im = _RAND_9619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9620 = {1{`RANDOM}};
  _T_5012_re = _RAND_9620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9621 = {1{`RANDOM}};
  _T_5012_im = _RAND_9621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9622 = {1{`RANDOM}};
  _T_5013_re = _RAND_9622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9623 = {1{`RANDOM}};
  _T_5013_im = _RAND_9623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9624 = {1{`RANDOM}};
  _T_5014_re = _RAND_9624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9625 = {1{`RANDOM}};
  _T_5014_im = _RAND_9625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9626 = {1{`RANDOM}};
  _T_5015_re = _RAND_9626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9627 = {1{`RANDOM}};
  _T_5015_im = _RAND_9627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9628 = {1{`RANDOM}};
  _T_5016_re = _RAND_9628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9629 = {1{`RANDOM}};
  _T_5016_im = _RAND_9629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9630 = {1{`RANDOM}};
  _T_5017_re = _RAND_9630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9631 = {1{`RANDOM}};
  _T_5017_im = _RAND_9631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9632 = {1{`RANDOM}};
  _T_5018_re = _RAND_9632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9633 = {1{`RANDOM}};
  _T_5018_im = _RAND_9633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9634 = {1{`RANDOM}};
  _T_5019_re = _RAND_9634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9635 = {1{`RANDOM}};
  _T_5019_im = _RAND_9635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9636 = {1{`RANDOM}};
  _T_5020_re = _RAND_9636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9637 = {1{`RANDOM}};
  _T_5020_im = _RAND_9637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9638 = {1{`RANDOM}};
  _T_5021_re = _RAND_9638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9639 = {1{`RANDOM}};
  _T_5021_im = _RAND_9639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9640 = {1{`RANDOM}};
  _T_5022_re = _RAND_9640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9641 = {1{`RANDOM}};
  _T_5022_im = _RAND_9641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9642 = {1{`RANDOM}};
  _T_5023_re = _RAND_9642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9643 = {1{`RANDOM}};
  _T_5023_im = _RAND_9643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9644 = {1{`RANDOM}};
  _T_5024_re = _RAND_9644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9645 = {1{`RANDOM}};
  _T_5024_im = _RAND_9645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9646 = {1{`RANDOM}};
  _T_5025_re = _RAND_9646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9647 = {1{`RANDOM}};
  _T_5025_im = _RAND_9647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9648 = {1{`RANDOM}};
  _T_5026_re = _RAND_9648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9649 = {1{`RANDOM}};
  _T_5026_im = _RAND_9649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9650 = {1{`RANDOM}};
  _T_5027_re = _RAND_9650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9651 = {1{`RANDOM}};
  _T_5027_im = _RAND_9651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9652 = {1{`RANDOM}};
  _T_5028_re = _RAND_9652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9653 = {1{`RANDOM}};
  _T_5028_im = _RAND_9653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9654 = {1{`RANDOM}};
  _T_5029_re = _RAND_9654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9655 = {1{`RANDOM}};
  _T_5029_im = _RAND_9655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9656 = {1{`RANDOM}};
  _T_5030_re = _RAND_9656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9657 = {1{`RANDOM}};
  _T_5030_im = _RAND_9657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9658 = {1{`RANDOM}};
  _T_5031_re = _RAND_9658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9659 = {1{`RANDOM}};
  _T_5031_im = _RAND_9659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9660 = {1{`RANDOM}};
  _T_5032_re = _RAND_9660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9661 = {1{`RANDOM}};
  _T_5032_im = _RAND_9661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9662 = {1{`RANDOM}};
  _T_5033_re = _RAND_9662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9663 = {1{`RANDOM}};
  _T_5033_im = _RAND_9663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9664 = {1{`RANDOM}};
  _T_5034_re = _RAND_9664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9665 = {1{`RANDOM}};
  _T_5034_im = _RAND_9665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9666 = {1{`RANDOM}};
  _T_5035_re = _RAND_9666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9667 = {1{`RANDOM}};
  _T_5035_im = _RAND_9667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9668 = {1{`RANDOM}};
  _T_5036_re = _RAND_9668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9669 = {1{`RANDOM}};
  _T_5036_im = _RAND_9669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9670 = {1{`RANDOM}};
  _T_5037_re = _RAND_9670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9671 = {1{`RANDOM}};
  _T_5037_im = _RAND_9671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9672 = {1{`RANDOM}};
  _T_5038_re = _RAND_9672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9673 = {1{`RANDOM}};
  _T_5038_im = _RAND_9673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9674 = {1{`RANDOM}};
  _T_5039_re = _RAND_9674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9675 = {1{`RANDOM}};
  _T_5039_im = _RAND_9675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9676 = {1{`RANDOM}};
  _T_5040_re = _RAND_9676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9677 = {1{`RANDOM}};
  _T_5040_im = _RAND_9677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9678 = {1{`RANDOM}};
  _T_5041_re = _RAND_9678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9679 = {1{`RANDOM}};
  _T_5041_im = _RAND_9679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9680 = {1{`RANDOM}};
  _T_5042_re = _RAND_9680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9681 = {1{`RANDOM}};
  _T_5042_im = _RAND_9681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9682 = {1{`RANDOM}};
  _T_5043_re = _RAND_9682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9683 = {1{`RANDOM}};
  _T_5043_im = _RAND_9683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9684 = {1{`RANDOM}};
  _T_5044_re = _RAND_9684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9685 = {1{`RANDOM}};
  _T_5044_im = _RAND_9685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9686 = {1{`RANDOM}};
  _T_5045_re = _RAND_9686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9687 = {1{`RANDOM}};
  _T_5045_im = _RAND_9687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9688 = {1{`RANDOM}};
  _T_5046_re = _RAND_9688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9689 = {1{`RANDOM}};
  _T_5046_im = _RAND_9689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9690 = {1{`RANDOM}};
  _T_5047_re = _RAND_9690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9691 = {1{`RANDOM}};
  _T_5047_im = _RAND_9691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9692 = {1{`RANDOM}};
  _T_5048_re = _RAND_9692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9693 = {1{`RANDOM}};
  _T_5048_im = _RAND_9693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9694 = {1{`RANDOM}};
  _T_5049_re = _RAND_9694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9695 = {1{`RANDOM}};
  _T_5049_im = _RAND_9695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9696 = {1{`RANDOM}};
  _T_5050_re = _RAND_9696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9697 = {1{`RANDOM}};
  _T_5050_im = _RAND_9697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9698 = {1{`RANDOM}};
  _T_5051_re = _RAND_9698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9699 = {1{`RANDOM}};
  _T_5051_im = _RAND_9699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9700 = {1{`RANDOM}};
  _T_5052_re = _RAND_9700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9701 = {1{`RANDOM}};
  _T_5052_im = _RAND_9701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9702 = {1{`RANDOM}};
  _T_5053_re = _RAND_9702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9703 = {1{`RANDOM}};
  _T_5053_im = _RAND_9703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9704 = {1{`RANDOM}};
  _T_5054_re = _RAND_9704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9705 = {1{`RANDOM}};
  _T_5054_im = _RAND_9705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9706 = {1{`RANDOM}};
  _T_5055_re = _RAND_9706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9707 = {1{`RANDOM}};
  _T_5055_im = _RAND_9707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9708 = {1{`RANDOM}};
  _T_5056_re = _RAND_9708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9709 = {1{`RANDOM}};
  _T_5056_im = _RAND_9709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9710 = {1{`RANDOM}};
  _T_5057_re = _RAND_9710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9711 = {1{`RANDOM}};
  _T_5057_im = _RAND_9711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9712 = {1{`RANDOM}};
  _T_5058_re = _RAND_9712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9713 = {1{`RANDOM}};
  _T_5058_im = _RAND_9713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9714 = {1{`RANDOM}};
  _T_5059_re = _RAND_9714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9715 = {1{`RANDOM}};
  _T_5059_im = _RAND_9715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9716 = {1{`RANDOM}};
  _T_5060_re = _RAND_9716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9717 = {1{`RANDOM}};
  _T_5060_im = _RAND_9717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9718 = {1{`RANDOM}};
  _T_5061_re = _RAND_9718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9719 = {1{`RANDOM}};
  _T_5061_im = _RAND_9719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9720 = {1{`RANDOM}};
  _T_5062_re = _RAND_9720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9721 = {1{`RANDOM}};
  _T_5062_im = _RAND_9721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9722 = {1{`RANDOM}};
  _T_5063_re = _RAND_9722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9723 = {1{`RANDOM}};
  _T_5063_im = _RAND_9723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9724 = {1{`RANDOM}};
  _T_5064_re = _RAND_9724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9725 = {1{`RANDOM}};
  _T_5064_im = _RAND_9725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9726 = {1{`RANDOM}};
  _T_5065_re = _RAND_9726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9727 = {1{`RANDOM}};
  _T_5065_im = _RAND_9727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9728 = {1{`RANDOM}};
  _T_5066_re = _RAND_9728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9729 = {1{`RANDOM}};
  _T_5066_im = _RAND_9729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9730 = {1{`RANDOM}};
  _T_5067_re = _RAND_9730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9731 = {1{`RANDOM}};
  _T_5067_im = _RAND_9731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9732 = {1{`RANDOM}};
  _T_5068_re = _RAND_9732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9733 = {1{`RANDOM}};
  _T_5068_im = _RAND_9733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9734 = {1{`RANDOM}};
  _T_5069_re = _RAND_9734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9735 = {1{`RANDOM}};
  _T_5069_im = _RAND_9735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9736 = {1{`RANDOM}};
  _T_5070_re = _RAND_9736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9737 = {1{`RANDOM}};
  _T_5070_im = _RAND_9737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9738 = {1{`RANDOM}};
  _T_5071_re = _RAND_9738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9739 = {1{`RANDOM}};
  _T_5071_im = _RAND_9739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9740 = {1{`RANDOM}};
  _T_5072_re = _RAND_9740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9741 = {1{`RANDOM}};
  _T_5072_im = _RAND_9741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9742 = {1{`RANDOM}};
  _T_5073_re = _RAND_9742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9743 = {1{`RANDOM}};
  _T_5073_im = _RAND_9743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9744 = {1{`RANDOM}};
  _T_5074_re = _RAND_9744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9745 = {1{`RANDOM}};
  _T_5074_im = _RAND_9745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9746 = {1{`RANDOM}};
  _T_5075_re = _RAND_9746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9747 = {1{`RANDOM}};
  _T_5075_im = _RAND_9747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9748 = {1{`RANDOM}};
  _T_5076_re = _RAND_9748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9749 = {1{`RANDOM}};
  _T_5076_im = _RAND_9749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9750 = {1{`RANDOM}};
  _T_5077_re = _RAND_9750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9751 = {1{`RANDOM}};
  _T_5077_im = _RAND_9751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9752 = {1{`RANDOM}};
  _T_5078_re = _RAND_9752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9753 = {1{`RANDOM}};
  _T_5078_im = _RAND_9753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9754 = {1{`RANDOM}};
  _T_5079_re = _RAND_9754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9755 = {1{`RANDOM}};
  _T_5079_im = _RAND_9755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9756 = {1{`RANDOM}};
  _T_5080_re = _RAND_9756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9757 = {1{`RANDOM}};
  _T_5080_im = _RAND_9757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9758 = {1{`RANDOM}};
  _T_5081_re = _RAND_9758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9759 = {1{`RANDOM}};
  _T_5081_im = _RAND_9759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9760 = {1{`RANDOM}};
  _T_5082_re = _RAND_9760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9761 = {1{`RANDOM}};
  _T_5082_im = _RAND_9761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9762 = {1{`RANDOM}};
  _T_5083_re = _RAND_9762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9763 = {1{`RANDOM}};
  _T_5083_im = _RAND_9763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9764 = {1{`RANDOM}};
  _T_5084_re = _RAND_9764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9765 = {1{`RANDOM}};
  _T_5084_im = _RAND_9765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9766 = {1{`RANDOM}};
  _T_5085_re = _RAND_9766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9767 = {1{`RANDOM}};
  _T_5085_im = _RAND_9767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9768 = {1{`RANDOM}};
  _T_5086_re = _RAND_9768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9769 = {1{`RANDOM}};
  _T_5086_im = _RAND_9769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9770 = {1{`RANDOM}};
  _T_5087_re = _RAND_9770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9771 = {1{`RANDOM}};
  _T_5087_im = _RAND_9771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9772 = {1{`RANDOM}};
  _T_5088_re = _RAND_9772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9773 = {1{`RANDOM}};
  _T_5088_im = _RAND_9773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9774 = {1{`RANDOM}};
  _T_5089_re = _RAND_9774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9775 = {1{`RANDOM}};
  _T_5089_im = _RAND_9775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9776 = {1{`RANDOM}};
  _T_5090_re = _RAND_9776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9777 = {1{`RANDOM}};
  _T_5090_im = _RAND_9777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9778 = {1{`RANDOM}};
  _T_5091_re = _RAND_9778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9779 = {1{`RANDOM}};
  _T_5091_im = _RAND_9779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9780 = {1{`RANDOM}};
  _T_5092_re = _RAND_9780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9781 = {1{`RANDOM}};
  _T_5092_im = _RAND_9781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9782 = {1{`RANDOM}};
  _T_5093_re = _RAND_9782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9783 = {1{`RANDOM}};
  _T_5093_im = _RAND_9783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9784 = {1{`RANDOM}};
  _T_5094_re = _RAND_9784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9785 = {1{`RANDOM}};
  _T_5094_im = _RAND_9785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9786 = {1{`RANDOM}};
  _T_5095_re = _RAND_9786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9787 = {1{`RANDOM}};
  _T_5095_im = _RAND_9787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9788 = {1{`RANDOM}};
  _T_5096_re = _RAND_9788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9789 = {1{`RANDOM}};
  _T_5096_im = _RAND_9789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9790 = {1{`RANDOM}};
  _T_5097_re = _RAND_9790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9791 = {1{`RANDOM}};
  _T_5097_im = _RAND_9791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9792 = {1{`RANDOM}};
  _T_5098_re = _RAND_9792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9793 = {1{`RANDOM}};
  _T_5098_im = _RAND_9793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9794 = {1{`RANDOM}};
  _T_5099_re = _RAND_9794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9795 = {1{`RANDOM}};
  _T_5099_im = _RAND_9795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9796 = {1{`RANDOM}};
  _T_5100_re = _RAND_9796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9797 = {1{`RANDOM}};
  _T_5100_im = _RAND_9797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9798 = {1{`RANDOM}};
  _T_5101_re = _RAND_9798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9799 = {1{`RANDOM}};
  _T_5101_im = _RAND_9799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9800 = {1{`RANDOM}};
  _T_5102_re = _RAND_9800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9801 = {1{`RANDOM}};
  _T_5102_im = _RAND_9801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9802 = {1{`RANDOM}};
  _T_5103_re = _RAND_9802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9803 = {1{`RANDOM}};
  _T_5103_im = _RAND_9803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9804 = {1{`RANDOM}};
  _T_5104_re = _RAND_9804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9805 = {1{`RANDOM}};
  _T_5104_im = _RAND_9805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9806 = {1{`RANDOM}};
  _T_5105_re = _RAND_9806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9807 = {1{`RANDOM}};
  _T_5105_im = _RAND_9807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9808 = {1{`RANDOM}};
  _T_5106_re = _RAND_9808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9809 = {1{`RANDOM}};
  _T_5106_im = _RAND_9809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9810 = {1{`RANDOM}};
  _T_5107_re = _RAND_9810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9811 = {1{`RANDOM}};
  _T_5107_im = _RAND_9811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9812 = {1{`RANDOM}};
  _T_5108_re = _RAND_9812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9813 = {1{`RANDOM}};
  _T_5108_im = _RAND_9813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9814 = {1{`RANDOM}};
  _T_5109_re = _RAND_9814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9815 = {1{`RANDOM}};
  _T_5109_im = _RAND_9815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9816 = {1{`RANDOM}};
  _T_5110_re = _RAND_9816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9817 = {1{`RANDOM}};
  _T_5110_im = _RAND_9817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9818 = {1{`RANDOM}};
  _T_5111_re = _RAND_9818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9819 = {1{`RANDOM}};
  _T_5111_im = _RAND_9819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9820 = {1{`RANDOM}};
  _T_5112_re = _RAND_9820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9821 = {1{`RANDOM}};
  _T_5112_im = _RAND_9821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9822 = {1{`RANDOM}};
  _T_5113_re = _RAND_9822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9823 = {1{`RANDOM}};
  _T_5113_im = _RAND_9823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9824 = {1{`RANDOM}};
  _T_5114_re = _RAND_9824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9825 = {1{`RANDOM}};
  _T_5114_im = _RAND_9825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9826 = {1{`RANDOM}};
  _T_5115_re = _RAND_9826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9827 = {1{`RANDOM}};
  _T_5115_im = _RAND_9827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9828 = {1{`RANDOM}};
  _T_5116_re = _RAND_9828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9829 = {1{`RANDOM}};
  _T_5116_im = _RAND_9829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9830 = {1{`RANDOM}};
  _T_5117_re = _RAND_9830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9831 = {1{`RANDOM}};
  _T_5117_im = _RAND_9831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9832 = {1{`RANDOM}};
  _T_5118_re = _RAND_9832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9833 = {1{`RANDOM}};
  _T_5118_im = _RAND_9833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9834 = {1{`RANDOM}};
  _T_5119_re = _RAND_9834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9835 = {1{`RANDOM}};
  _T_5119_im = _RAND_9835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9836 = {1{`RANDOM}};
  _T_5120_re = _RAND_9836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9837 = {1{`RANDOM}};
  _T_5120_im = _RAND_9837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9838 = {1{`RANDOM}};
  _T_5121_re = _RAND_9838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9839 = {1{`RANDOM}};
  _T_5121_im = _RAND_9839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9840 = {1{`RANDOM}};
  _T_5122_re = _RAND_9840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9841 = {1{`RANDOM}};
  _T_5122_im = _RAND_9841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9842 = {1{`RANDOM}};
  _T_5123_re = _RAND_9842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9843 = {1{`RANDOM}};
  _T_5123_im = _RAND_9843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9844 = {1{`RANDOM}};
  _T_5124_re = _RAND_9844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9845 = {1{`RANDOM}};
  _T_5124_im = _RAND_9845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9846 = {1{`RANDOM}};
  _T_5125_re = _RAND_9846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9847 = {1{`RANDOM}};
  _T_5125_im = _RAND_9847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9848 = {1{`RANDOM}};
  _T_5126_re = _RAND_9848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9849 = {1{`RANDOM}};
  _T_5126_im = _RAND_9849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9850 = {1{`RANDOM}};
  _T_5127_re = _RAND_9850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9851 = {1{`RANDOM}};
  _T_5127_im = _RAND_9851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9852 = {1{`RANDOM}};
  _T_5128_re = _RAND_9852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9853 = {1{`RANDOM}};
  _T_5128_im = _RAND_9853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9854 = {1{`RANDOM}};
  _T_5129_re = _RAND_9854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9855 = {1{`RANDOM}};
  _T_5129_im = _RAND_9855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9856 = {1{`RANDOM}};
  _T_5130_re = _RAND_9856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9857 = {1{`RANDOM}};
  _T_5130_im = _RAND_9857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9858 = {1{`RANDOM}};
  _T_5131_re = _RAND_9858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9859 = {1{`RANDOM}};
  _T_5131_im = _RAND_9859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9860 = {1{`RANDOM}};
  _T_5132_re = _RAND_9860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9861 = {1{`RANDOM}};
  _T_5132_im = _RAND_9861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9862 = {1{`RANDOM}};
  _T_5133_re = _RAND_9862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9863 = {1{`RANDOM}};
  _T_5133_im = _RAND_9863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9864 = {1{`RANDOM}};
  _T_5134_re = _RAND_9864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9865 = {1{`RANDOM}};
  _T_5134_im = _RAND_9865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9866 = {1{`RANDOM}};
  _T_5135_re = _RAND_9866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9867 = {1{`RANDOM}};
  _T_5135_im = _RAND_9867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9868 = {1{`RANDOM}};
  _T_5136_re = _RAND_9868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9869 = {1{`RANDOM}};
  _T_5136_im = _RAND_9869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9870 = {1{`RANDOM}};
  _T_5137_re = _RAND_9870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9871 = {1{`RANDOM}};
  _T_5137_im = _RAND_9871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9872 = {1{`RANDOM}};
  _T_5138_re = _RAND_9872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9873 = {1{`RANDOM}};
  _T_5138_im = _RAND_9873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9874 = {1{`RANDOM}};
  _T_5139_re = _RAND_9874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9875 = {1{`RANDOM}};
  _T_5139_im = _RAND_9875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9876 = {1{`RANDOM}};
  _T_5140_re = _RAND_9876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9877 = {1{`RANDOM}};
  _T_5140_im = _RAND_9877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9878 = {1{`RANDOM}};
  _T_5141_re = _RAND_9878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9879 = {1{`RANDOM}};
  _T_5141_im = _RAND_9879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9880 = {1{`RANDOM}};
  _T_5142_re = _RAND_9880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9881 = {1{`RANDOM}};
  _T_5142_im = _RAND_9881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9882 = {1{`RANDOM}};
  _T_5143_re = _RAND_9882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9883 = {1{`RANDOM}};
  _T_5143_im = _RAND_9883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9884 = {1{`RANDOM}};
  _T_5144_re = _RAND_9884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9885 = {1{`RANDOM}};
  _T_5144_im = _RAND_9885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9886 = {1{`RANDOM}};
  _T_5145_re = _RAND_9886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9887 = {1{`RANDOM}};
  _T_5145_im = _RAND_9887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9888 = {1{`RANDOM}};
  _T_5146_re = _RAND_9888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9889 = {1{`RANDOM}};
  _T_5146_im = _RAND_9889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9890 = {1{`RANDOM}};
  _T_5147_re = _RAND_9890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9891 = {1{`RANDOM}};
  _T_5147_im = _RAND_9891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9892 = {1{`RANDOM}};
  _T_5148_re = _RAND_9892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9893 = {1{`RANDOM}};
  _T_5148_im = _RAND_9893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9894 = {1{`RANDOM}};
  _T_5149_re = _RAND_9894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9895 = {1{`RANDOM}};
  _T_5149_im = _RAND_9895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9896 = {1{`RANDOM}};
  _T_5150_re = _RAND_9896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9897 = {1{`RANDOM}};
  _T_5150_im = _RAND_9897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9898 = {1{`RANDOM}};
  _T_5151_re = _RAND_9898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9899 = {1{`RANDOM}};
  _T_5151_im = _RAND_9899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9900 = {1{`RANDOM}};
  _T_5152_re = _RAND_9900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9901 = {1{`RANDOM}};
  _T_5152_im = _RAND_9901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9902 = {1{`RANDOM}};
  _T_5153_re = _RAND_9902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9903 = {1{`RANDOM}};
  _T_5153_im = _RAND_9903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9904 = {1{`RANDOM}};
  _T_5154_re = _RAND_9904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9905 = {1{`RANDOM}};
  _T_5154_im = _RAND_9905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9906 = {1{`RANDOM}};
  _T_5155_re = _RAND_9906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9907 = {1{`RANDOM}};
  _T_5155_im = _RAND_9907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9908 = {1{`RANDOM}};
  _T_5156_re = _RAND_9908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9909 = {1{`RANDOM}};
  _T_5156_im = _RAND_9909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9910 = {1{`RANDOM}};
  _T_5157_re = _RAND_9910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9911 = {1{`RANDOM}};
  _T_5157_im = _RAND_9911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9912 = {1{`RANDOM}};
  _T_5158_re = _RAND_9912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9913 = {1{`RANDOM}};
  _T_5158_im = _RAND_9913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9914 = {1{`RANDOM}};
  _T_5159_re = _RAND_9914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9915 = {1{`RANDOM}};
  _T_5159_im = _RAND_9915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9916 = {1{`RANDOM}};
  _T_5160_re = _RAND_9916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9917 = {1{`RANDOM}};
  _T_5160_im = _RAND_9917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9918 = {1{`RANDOM}};
  _T_5161_re = _RAND_9918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9919 = {1{`RANDOM}};
  _T_5161_im = _RAND_9919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9920 = {1{`RANDOM}};
  _T_5162_re = _RAND_9920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9921 = {1{`RANDOM}};
  _T_5162_im = _RAND_9921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9922 = {1{`RANDOM}};
  _T_5163_re = _RAND_9922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9923 = {1{`RANDOM}};
  _T_5163_im = _RAND_9923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9924 = {1{`RANDOM}};
  _T_5164_re = _RAND_9924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9925 = {1{`RANDOM}};
  _T_5164_im = _RAND_9925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9926 = {1{`RANDOM}};
  _T_5165_re = _RAND_9926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9927 = {1{`RANDOM}};
  _T_5165_im = _RAND_9927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9928 = {1{`RANDOM}};
  _T_5166_re = _RAND_9928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9929 = {1{`RANDOM}};
  _T_5166_im = _RAND_9929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9930 = {1{`RANDOM}};
  _T_5167_re = _RAND_9930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9931 = {1{`RANDOM}};
  _T_5167_im = _RAND_9931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9932 = {1{`RANDOM}};
  _T_5168_re = _RAND_9932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9933 = {1{`RANDOM}};
  _T_5168_im = _RAND_9933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9934 = {1{`RANDOM}};
  _T_5169_re = _RAND_9934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9935 = {1{`RANDOM}};
  _T_5169_im = _RAND_9935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9936 = {1{`RANDOM}};
  _T_5170_re = _RAND_9936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9937 = {1{`RANDOM}};
  _T_5170_im = _RAND_9937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9938 = {1{`RANDOM}};
  _T_5171_re = _RAND_9938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9939 = {1{`RANDOM}};
  _T_5171_im = _RAND_9939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9940 = {1{`RANDOM}};
  _T_5172_re = _RAND_9940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9941 = {1{`RANDOM}};
  _T_5172_im = _RAND_9941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9942 = {1{`RANDOM}};
  _T_5173_re = _RAND_9942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9943 = {1{`RANDOM}};
  _T_5173_im = _RAND_9943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9944 = {1{`RANDOM}};
  _T_5174_re = _RAND_9944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9945 = {1{`RANDOM}};
  _T_5174_im = _RAND_9945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9946 = {1{`RANDOM}};
  _T_5175_re = _RAND_9946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9947 = {1{`RANDOM}};
  _T_5175_im = _RAND_9947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9948 = {1{`RANDOM}};
  _T_5176_re = _RAND_9948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9949 = {1{`RANDOM}};
  _T_5176_im = _RAND_9949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9950 = {1{`RANDOM}};
  _T_5177_re = _RAND_9950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9951 = {1{`RANDOM}};
  _T_5177_im = _RAND_9951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9952 = {1{`RANDOM}};
  _T_5178_re = _RAND_9952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9953 = {1{`RANDOM}};
  _T_5178_im = _RAND_9953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9954 = {1{`RANDOM}};
  _T_5179_re = _RAND_9954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9955 = {1{`RANDOM}};
  _T_5179_im = _RAND_9955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9956 = {1{`RANDOM}};
  _T_5180_re = _RAND_9956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9957 = {1{`RANDOM}};
  _T_5180_im = _RAND_9957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9958 = {1{`RANDOM}};
  _T_5181_re = _RAND_9958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9959 = {1{`RANDOM}};
  _T_5181_im = _RAND_9959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9960 = {1{`RANDOM}};
  _T_5182_re = _RAND_9960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9961 = {1{`RANDOM}};
  _T_5182_im = _RAND_9961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9962 = {1{`RANDOM}};
  _T_5183_re = _RAND_9962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9963 = {1{`RANDOM}};
  _T_5183_im = _RAND_9963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9964 = {1{`RANDOM}};
  _T_5184_re = _RAND_9964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9965 = {1{`RANDOM}};
  _T_5184_im = _RAND_9965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9966 = {1{`RANDOM}};
  _T_5185_re = _RAND_9966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9967 = {1{`RANDOM}};
  _T_5185_im = _RAND_9967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9968 = {1{`RANDOM}};
  _T_5186_re = _RAND_9968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9969 = {1{`RANDOM}};
  _T_5186_im = _RAND_9969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9970 = {1{`RANDOM}};
  _T_5187_re = _RAND_9970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9971 = {1{`RANDOM}};
  _T_5187_im = _RAND_9971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9972 = {1{`RANDOM}};
  _T_5188_re = _RAND_9972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9973 = {1{`RANDOM}};
  _T_5188_im = _RAND_9973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9974 = {1{`RANDOM}};
  _T_5189_re = _RAND_9974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9975 = {1{`RANDOM}};
  _T_5189_im = _RAND_9975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9976 = {1{`RANDOM}};
  _T_5190_re = _RAND_9976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9977 = {1{`RANDOM}};
  _T_5190_im = _RAND_9977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9978 = {1{`RANDOM}};
  _T_5191_re = _RAND_9978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9979 = {1{`RANDOM}};
  _T_5191_im = _RAND_9979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9980 = {1{`RANDOM}};
  _T_5192_re = _RAND_9980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9981 = {1{`RANDOM}};
  _T_5192_im = _RAND_9981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9982 = {1{`RANDOM}};
  _T_5193_re = _RAND_9982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9983 = {1{`RANDOM}};
  _T_5193_im = _RAND_9983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9984 = {1{`RANDOM}};
  _T_5194_re = _RAND_9984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9985 = {1{`RANDOM}};
  _T_5194_im = _RAND_9985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9986 = {1{`RANDOM}};
  _T_5195_re = _RAND_9986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9987 = {1{`RANDOM}};
  _T_5195_im = _RAND_9987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9988 = {1{`RANDOM}};
  _T_5196_re = _RAND_9988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9989 = {1{`RANDOM}};
  _T_5196_im = _RAND_9989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9990 = {1{`RANDOM}};
  _T_5197_re = _RAND_9990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9991 = {1{`RANDOM}};
  _T_5197_im = _RAND_9991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9992 = {1{`RANDOM}};
  _T_5198_re = _RAND_9992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9993 = {1{`RANDOM}};
  _T_5198_im = _RAND_9993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9994 = {1{`RANDOM}};
  _T_5199_re = _RAND_9994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9995 = {1{`RANDOM}};
  _T_5199_im = _RAND_9995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9996 = {1{`RANDOM}};
  _T_5200_re = _RAND_9996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9997 = {1{`RANDOM}};
  _T_5200_im = _RAND_9997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9998 = {1{`RANDOM}};
  _T_5201_re = _RAND_9998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9999 = {1{`RANDOM}};
  _T_5201_im = _RAND_9999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10000 = {1{`RANDOM}};
  _T_5202_re = _RAND_10000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10001 = {1{`RANDOM}};
  _T_5202_im = _RAND_10001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10002 = {1{`RANDOM}};
  _T_5203_re = _RAND_10002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10003 = {1{`RANDOM}};
  _T_5203_im = _RAND_10003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10004 = {1{`RANDOM}};
  _T_5204_re = _RAND_10004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10005 = {1{`RANDOM}};
  _T_5204_im = _RAND_10005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10006 = {1{`RANDOM}};
  _T_5205_re = _RAND_10006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10007 = {1{`RANDOM}};
  _T_5205_im = _RAND_10007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10008 = {1{`RANDOM}};
  _T_5206_re = _RAND_10008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10009 = {1{`RANDOM}};
  _T_5206_im = _RAND_10009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10010 = {1{`RANDOM}};
  _T_5207_re = _RAND_10010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10011 = {1{`RANDOM}};
  _T_5207_im = _RAND_10011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10012 = {1{`RANDOM}};
  _T_5208_re = _RAND_10012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10013 = {1{`RANDOM}};
  _T_5208_im = _RAND_10013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10014 = {1{`RANDOM}};
  _T_5209_re = _RAND_10014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10015 = {1{`RANDOM}};
  _T_5209_im = _RAND_10015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10016 = {1{`RANDOM}};
  _T_5210_re = _RAND_10016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10017 = {1{`RANDOM}};
  _T_5210_im = _RAND_10017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10018 = {1{`RANDOM}};
  _T_5211_re = _RAND_10018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10019 = {1{`RANDOM}};
  _T_5211_im = _RAND_10019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10020 = {1{`RANDOM}};
  _T_5212_re = _RAND_10020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10021 = {1{`RANDOM}};
  _T_5212_im = _RAND_10021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10022 = {1{`RANDOM}};
  _T_5213_re = _RAND_10022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10023 = {1{`RANDOM}};
  _T_5213_im = _RAND_10023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10024 = {1{`RANDOM}};
  _T_5214_re = _RAND_10024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10025 = {1{`RANDOM}};
  _T_5214_im = _RAND_10025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10026 = {1{`RANDOM}};
  _T_5215_re = _RAND_10026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10027 = {1{`RANDOM}};
  _T_5215_im = _RAND_10027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10028 = {1{`RANDOM}};
  _T_5216_re = _RAND_10028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10029 = {1{`RANDOM}};
  _T_5216_im = _RAND_10029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10030 = {1{`RANDOM}};
  _T_5217_re = _RAND_10030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10031 = {1{`RANDOM}};
  _T_5217_im = _RAND_10031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10032 = {1{`RANDOM}};
  _T_5218_re = _RAND_10032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10033 = {1{`RANDOM}};
  _T_5218_im = _RAND_10033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10034 = {1{`RANDOM}};
  _T_5219_re = _RAND_10034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10035 = {1{`RANDOM}};
  _T_5219_im = _RAND_10035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10036 = {1{`RANDOM}};
  _T_5220_re = _RAND_10036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10037 = {1{`RANDOM}};
  _T_5220_im = _RAND_10037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10038 = {1{`RANDOM}};
  _T_5221_re = _RAND_10038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10039 = {1{`RANDOM}};
  _T_5221_im = _RAND_10039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10040 = {1{`RANDOM}};
  _T_5222_re = _RAND_10040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10041 = {1{`RANDOM}};
  _T_5222_im = _RAND_10041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10042 = {1{`RANDOM}};
  _T_5223_re = _RAND_10042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10043 = {1{`RANDOM}};
  _T_5223_im = _RAND_10043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10044 = {1{`RANDOM}};
  _T_5224_re = _RAND_10044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10045 = {1{`RANDOM}};
  _T_5224_im = _RAND_10045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10046 = {1{`RANDOM}};
  _T_5225_re = _RAND_10046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10047 = {1{`RANDOM}};
  _T_5225_im = _RAND_10047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10048 = {1{`RANDOM}};
  _T_5226_re = _RAND_10048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10049 = {1{`RANDOM}};
  _T_5226_im = _RAND_10049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10050 = {1{`RANDOM}};
  _T_5227_re = _RAND_10050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10051 = {1{`RANDOM}};
  _T_5227_im = _RAND_10051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10052 = {1{`RANDOM}};
  _T_5228_re = _RAND_10052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10053 = {1{`RANDOM}};
  _T_5228_im = _RAND_10053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10054 = {1{`RANDOM}};
  _T_5229_re = _RAND_10054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10055 = {1{`RANDOM}};
  _T_5229_im = _RAND_10055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10056 = {1{`RANDOM}};
  _T_5230_re = _RAND_10056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10057 = {1{`RANDOM}};
  _T_5230_im = _RAND_10057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10058 = {1{`RANDOM}};
  _T_5231_re = _RAND_10058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10059 = {1{`RANDOM}};
  _T_5231_im = _RAND_10059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10060 = {1{`RANDOM}};
  _T_5232_re = _RAND_10060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10061 = {1{`RANDOM}};
  _T_5232_im = _RAND_10061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10062 = {1{`RANDOM}};
  _T_5233_re = _RAND_10062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10063 = {1{`RANDOM}};
  _T_5233_im = _RAND_10063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10064 = {1{`RANDOM}};
  _T_5234_re = _RAND_10064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10065 = {1{`RANDOM}};
  _T_5234_im = _RAND_10065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10066 = {1{`RANDOM}};
  _T_5235_re = _RAND_10066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10067 = {1{`RANDOM}};
  _T_5235_im = _RAND_10067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10068 = {1{`RANDOM}};
  _T_5236_re = _RAND_10068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10069 = {1{`RANDOM}};
  _T_5236_im = _RAND_10069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10070 = {1{`RANDOM}};
  _T_5237_re = _RAND_10070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10071 = {1{`RANDOM}};
  _T_5237_im = _RAND_10071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10072 = {1{`RANDOM}};
  _T_5238_re = _RAND_10072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10073 = {1{`RANDOM}};
  _T_5238_im = _RAND_10073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10074 = {1{`RANDOM}};
  _T_5239_re = _RAND_10074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10075 = {1{`RANDOM}};
  _T_5239_im = _RAND_10075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10076 = {1{`RANDOM}};
  _T_5240_re = _RAND_10076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10077 = {1{`RANDOM}};
  _T_5240_im = _RAND_10077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10078 = {1{`RANDOM}};
  _T_5241_re = _RAND_10078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10079 = {1{`RANDOM}};
  _T_5241_im = _RAND_10079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10080 = {1{`RANDOM}};
  _T_5242_re = _RAND_10080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10081 = {1{`RANDOM}};
  _T_5242_im = _RAND_10081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10082 = {1{`RANDOM}};
  _T_5243_re = _RAND_10082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10083 = {1{`RANDOM}};
  _T_5243_im = _RAND_10083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10084 = {1{`RANDOM}};
  _T_5244_re = _RAND_10084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10085 = {1{`RANDOM}};
  _T_5244_im = _RAND_10085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10086 = {1{`RANDOM}};
  _T_5245_re = _RAND_10086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10087 = {1{`RANDOM}};
  _T_5245_im = _RAND_10087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10088 = {1{`RANDOM}};
  _T_5246_re = _RAND_10088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10089 = {1{`RANDOM}};
  _T_5246_im = _RAND_10089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10090 = {1{`RANDOM}};
  _T_5247_re = _RAND_10090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10091 = {1{`RANDOM}};
  _T_5247_im = _RAND_10091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10092 = {1{`RANDOM}};
  _T_5248_re = _RAND_10092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10093 = {1{`RANDOM}};
  _T_5248_im = _RAND_10093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10094 = {1{`RANDOM}};
  _T_5249_re = _RAND_10094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10095 = {1{`RANDOM}};
  _T_5249_im = _RAND_10095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10096 = {1{`RANDOM}};
  _T_5250_re = _RAND_10096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10097 = {1{`RANDOM}};
  _T_5250_im = _RAND_10097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10098 = {1{`RANDOM}};
  _T_5251_re = _RAND_10098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10099 = {1{`RANDOM}};
  _T_5251_im = _RAND_10099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10100 = {1{`RANDOM}};
  _T_5252_re = _RAND_10100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10101 = {1{`RANDOM}};
  _T_5252_im = _RAND_10101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10102 = {1{`RANDOM}};
  _T_5253_re = _RAND_10102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10103 = {1{`RANDOM}};
  _T_5253_im = _RAND_10103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10104 = {1{`RANDOM}};
  _T_5254_re = _RAND_10104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10105 = {1{`RANDOM}};
  _T_5254_im = _RAND_10105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10106 = {1{`RANDOM}};
  _T_5255_re = _RAND_10106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10107 = {1{`RANDOM}};
  _T_5255_im = _RAND_10107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10108 = {1{`RANDOM}};
  _T_5256_re = _RAND_10108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10109 = {1{`RANDOM}};
  _T_5256_im = _RAND_10109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10110 = {1{`RANDOM}};
  _T_5257_re = _RAND_10110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10111 = {1{`RANDOM}};
  _T_5257_im = _RAND_10111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10112 = {1{`RANDOM}};
  _T_5258_re = _RAND_10112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10113 = {1{`RANDOM}};
  _T_5258_im = _RAND_10113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10114 = {1{`RANDOM}};
  _T_5259_re = _RAND_10114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10115 = {1{`RANDOM}};
  _T_5259_im = _RAND_10115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10116 = {1{`RANDOM}};
  _T_5260_re = _RAND_10116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10117 = {1{`RANDOM}};
  _T_5260_im = _RAND_10117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10118 = {1{`RANDOM}};
  _T_5261_re = _RAND_10118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10119 = {1{`RANDOM}};
  _T_5261_im = _RAND_10119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10120 = {1{`RANDOM}};
  _T_5262_re = _RAND_10120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10121 = {1{`RANDOM}};
  _T_5262_im = _RAND_10121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10122 = {1{`RANDOM}};
  _T_5263_re = _RAND_10122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10123 = {1{`RANDOM}};
  _T_5263_im = _RAND_10123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10124 = {1{`RANDOM}};
  _T_5264_re = _RAND_10124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10125 = {1{`RANDOM}};
  _T_5264_im = _RAND_10125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10126 = {1{`RANDOM}};
  _T_5265_re = _RAND_10126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10127 = {1{`RANDOM}};
  _T_5265_im = _RAND_10127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10128 = {1{`RANDOM}};
  _T_5266_re = _RAND_10128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10129 = {1{`RANDOM}};
  _T_5266_im = _RAND_10129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10130 = {1{`RANDOM}};
  _T_5267_re = _RAND_10130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10131 = {1{`RANDOM}};
  _T_5267_im = _RAND_10131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10132 = {1{`RANDOM}};
  _T_5268_re = _RAND_10132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10133 = {1{`RANDOM}};
  _T_5268_im = _RAND_10133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10134 = {1{`RANDOM}};
  _T_5269_re = _RAND_10134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10135 = {1{`RANDOM}};
  _T_5269_im = _RAND_10135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10136 = {1{`RANDOM}};
  _T_5270_re = _RAND_10136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10137 = {1{`RANDOM}};
  _T_5270_im = _RAND_10137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10138 = {1{`RANDOM}};
  _T_5271_re = _RAND_10138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10139 = {1{`RANDOM}};
  _T_5271_im = _RAND_10139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10140 = {1{`RANDOM}};
  _T_5272_re = _RAND_10140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10141 = {1{`RANDOM}};
  _T_5272_im = _RAND_10141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10142 = {1{`RANDOM}};
  _T_5273_re = _RAND_10142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10143 = {1{`RANDOM}};
  _T_5273_im = _RAND_10143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10144 = {1{`RANDOM}};
  _T_5274_re = _RAND_10144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10145 = {1{`RANDOM}};
  _T_5274_im = _RAND_10145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10146 = {1{`RANDOM}};
  _T_5275_re = _RAND_10146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10147 = {1{`RANDOM}};
  _T_5275_im = _RAND_10147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10148 = {1{`RANDOM}};
  _T_5276_re = _RAND_10148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10149 = {1{`RANDOM}};
  _T_5276_im = _RAND_10149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10150 = {1{`RANDOM}};
  _T_5277_re = _RAND_10150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10151 = {1{`RANDOM}};
  _T_5277_im = _RAND_10151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10152 = {1{`RANDOM}};
  _T_5278_re = _RAND_10152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10153 = {1{`RANDOM}};
  _T_5278_im = _RAND_10153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10154 = {1{`RANDOM}};
  _T_5279_re = _RAND_10154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10155 = {1{`RANDOM}};
  _T_5279_im = _RAND_10155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10156 = {1{`RANDOM}};
  _T_5280_re = _RAND_10156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10157 = {1{`RANDOM}};
  _T_5280_im = _RAND_10157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10158 = {1{`RANDOM}};
  _T_5281_re = _RAND_10158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10159 = {1{`RANDOM}};
  _T_5281_im = _RAND_10159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10160 = {1{`RANDOM}};
  _T_5282_re = _RAND_10160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10161 = {1{`RANDOM}};
  _T_5282_im = _RAND_10161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10162 = {1{`RANDOM}};
  _T_5283_re = _RAND_10162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10163 = {1{`RANDOM}};
  _T_5283_im = _RAND_10163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10164 = {1{`RANDOM}};
  _T_5284_re = _RAND_10164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10165 = {1{`RANDOM}};
  _T_5284_im = _RAND_10165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10166 = {1{`RANDOM}};
  _T_5285_re = _RAND_10166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10167 = {1{`RANDOM}};
  _T_5285_im = _RAND_10167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10168 = {1{`RANDOM}};
  _T_5286_re = _RAND_10168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10169 = {1{`RANDOM}};
  _T_5286_im = _RAND_10169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10170 = {1{`RANDOM}};
  _T_5287_re = _RAND_10170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10171 = {1{`RANDOM}};
  _T_5287_im = _RAND_10171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10172 = {1{`RANDOM}};
  _T_5288_re = _RAND_10172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10173 = {1{`RANDOM}};
  _T_5288_im = _RAND_10173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10174 = {1{`RANDOM}};
  _T_5289_re = _RAND_10174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10175 = {1{`RANDOM}};
  _T_5289_im = _RAND_10175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10176 = {1{`RANDOM}};
  _T_5290_re = _RAND_10176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10177 = {1{`RANDOM}};
  _T_5290_im = _RAND_10177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10178 = {1{`RANDOM}};
  _T_5291_re = _RAND_10178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10179 = {1{`RANDOM}};
  _T_5291_im = _RAND_10179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10180 = {1{`RANDOM}};
  _T_5292_re = _RAND_10180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10181 = {1{`RANDOM}};
  _T_5292_im = _RAND_10181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10182 = {1{`RANDOM}};
  _T_5293_re = _RAND_10182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10183 = {1{`RANDOM}};
  _T_5293_im = _RAND_10183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10184 = {1{`RANDOM}};
  _T_5294_re = _RAND_10184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10185 = {1{`RANDOM}};
  _T_5294_im = _RAND_10185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10186 = {1{`RANDOM}};
  _T_5295_re = _RAND_10186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10187 = {1{`RANDOM}};
  _T_5295_im = _RAND_10187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10188 = {1{`RANDOM}};
  _T_5296_re = _RAND_10188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10189 = {1{`RANDOM}};
  _T_5296_im = _RAND_10189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10190 = {1{`RANDOM}};
  _T_5297_re = _RAND_10190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10191 = {1{`RANDOM}};
  _T_5297_im = _RAND_10191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10192 = {1{`RANDOM}};
  _T_5298_re = _RAND_10192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10193 = {1{`RANDOM}};
  _T_5298_im = _RAND_10193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10194 = {1{`RANDOM}};
  _T_5299_re = _RAND_10194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10195 = {1{`RANDOM}};
  _T_5299_im = _RAND_10195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10196 = {1{`RANDOM}};
  _T_5300_re = _RAND_10196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10197 = {1{`RANDOM}};
  _T_5300_im = _RAND_10197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10198 = {1{`RANDOM}};
  _T_5301_re = _RAND_10198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10199 = {1{`RANDOM}};
  _T_5301_im = _RAND_10199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10200 = {1{`RANDOM}};
  _T_5302_re = _RAND_10200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10201 = {1{`RANDOM}};
  _T_5302_im = _RAND_10201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10202 = {1{`RANDOM}};
  _T_5303_re = _RAND_10202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10203 = {1{`RANDOM}};
  _T_5303_im = _RAND_10203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10204 = {1{`RANDOM}};
  _T_5304_re = _RAND_10204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10205 = {1{`RANDOM}};
  _T_5304_im = _RAND_10205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10206 = {1{`RANDOM}};
  _T_5305_re = _RAND_10206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10207 = {1{`RANDOM}};
  _T_5305_im = _RAND_10207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10208 = {1{`RANDOM}};
  _T_5306_re = _RAND_10208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10209 = {1{`RANDOM}};
  _T_5306_im = _RAND_10209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10210 = {1{`RANDOM}};
  _T_5307_re = _RAND_10210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10211 = {1{`RANDOM}};
  _T_5307_im = _RAND_10211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10212 = {1{`RANDOM}};
  _T_5308_re = _RAND_10212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10213 = {1{`RANDOM}};
  _T_5308_im = _RAND_10213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10214 = {1{`RANDOM}};
  _T_5309_re = _RAND_10214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10215 = {1{`RANDOM}};
  _T_5309_im = _RAND_10215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10216 = {1{`RANDOM}};
  _T_5310_re = _RAND_10216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10217 = {1{`RANDOM}};
  _T_5310_im = _RAND_10217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10218 = {1{`RANDOM}};
  _T_5311_re = _RAND_10218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10219 = {1{`RANDOM}};
  _T_5311_im = _RAND_10219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10220 = {1{`RANDOM}};
  _T_5312_re = _RAND_10220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10221 = {1{`RANDOM}};
  _T_5312_im = _RAND_10221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10222 = {1{`RANDOM}};
  _T_5313_re = _RAND_10222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10223 = {1{`RANDOM}};
  _T_5313_im = _RAND_10223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10224 = {1{`RANDOM}};
  _T_5314_re = _RAND_10224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10225 = {1{`RANDOM}};
  _T_5314_im = _RAND_10225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10226 = {1{`RANDOM}};
  _T_5315_re = _RAND_10226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10227 = {1{`RANDOM}};
  _T_5315_im = _RAND_10227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10228 = {1{`RANDOM}};
  _T_5316_re = _RAND_10228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10229 = {1{`RANDOM}};
  _T_5316_im = _RAND_10229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10230 = {1{`RANDOM}};
  _T_5317_re = _RAND_10230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10231 = {1{`RANDOM}};
  _T_5317_im = _RAND_10231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10232 = {1{`RANDOM}};
  _T_5318_re = _RAND_10232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10233 = {1{`RANDOM}};
  _T_5318_im = _RAND_10233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10234 = {1{`RANDOM}};
  _T_5319_re = _RAND_10234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10235 = {1{`RANDOM}};
  _T_5319_im = _RAND_10235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10236 = {1{`RANDOM}};
  _T_5320_re = _RAND_10236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10237 = {1{`RANDOM}};
  _T_5320_im = _RAND_10237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10238 = {1{`RANDOM}};
  _T_5321_re = _RAND_10238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10239 = {1{`RANDOM}};
  _T_5321_im = _RAND_10239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10240 = {1{`RANDOM}};
  _T_5322_re = _RAND_10240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10241 = {1{`RANDOM}};
  _T_5322_im = _RAND_10241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10242 = {1{`RANDOM}};
  _T_5325_re = _RAND_10242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10243 = {1{`RANDOM}};
  _T_5325_im = _RAND_10243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10244 = {1{`RANDOM}};
  _T_5326_re = _RAND_10244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10245 = {1{`RANDOM}};
  _T_5326_im = _RAND_10245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10246 = {1{`RANDOM}};
  _T_5327_re = _RAND_10246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10247 = {1{`RANDOM}};
  _T_5327_im = _RAND_10247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10248 = {1{`RANDOM}};
  _T_5328_re = _RAND_10248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10249 = {1{`RANDOM}};
  _T_5328_im = _RAND_10249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10250 = {1{`RANDOM}};
  _T_5329_re = _RAND_10250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10251 = {1{`RANDOM}};
  _T_5329_im = _RAND_10251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10252 = {1{`RANDOM}};
  _T_5330_re = _RAND_10252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10253 = {1{`RANDOM}};
  _T_5330_im = _RAND_10253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10254 = {1{`RANDOM}};
  _T_5331_re = _RAND_10254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10255 = {1{`RANDOM}};
  _T_5331_im = _RAND_10255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10256 = {1{`RANDOM}};
  _T_5332_re = _RAND_10256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10257 = {1{`RANDOM}};
  _T_5332_im = _RAND_10257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10258 = {1{`RANDOM}};
  _T_5333_re = _RAND_10258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10259 = {1{`RANDOM}};
  _T_5333_im = _RAND_10259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10260 = {1{`RANDOM}};
  _T_5334_re = _RAND_10260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10261 = {1{`RANDOM}};
  _T_5334_im = _RAND_10261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10262 = {1{`RANDOM}};
  _T_5335_re = _RAND_10262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10263 = {1{`RANDOM}};
  _T_5335_im = _RAND_10263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10264 = {1{`RANDOM}};
  _T_5336_re = _RAND_10264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10265 = {1{`RANDOM}};
  _T_5336_im = _RAND_10265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10266 = {1{`RANDOM}};
  _T_5337_re = _RAND_10266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10267 = {1{`RANDOM}};
  _T_5337_im = _RAND_10267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10268 = {1{`RANDOM}};
  _T_5338_re = _RAND_10268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10269 = {1{`RANDOM}};
  _T_5338_im = _RAND_10269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10270 = {1{`RANDOM}};
  _T_5339_re = _RAND_10270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10271 = {1{`RANDOM}};
  _T_5339_im = _RAND_10271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10272 = {1{`RANDOM}};
  _T_5340_re = _RAND_10272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10273 = {1{`RANDOM}};
  _T_5340_im = _RAND_10273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10274 = {1{`RANDOM}};
  _T_5341_re = _RAND_10274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10275 = {1{`RANDOM}};
  _T_5341_im = _RAND_10275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10276 = {1{`RANDOM}};
  _T_5342_re = _RAND_10276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10277 = {1{`RANDOM}};
  _T_5342_im = _RAND_10277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10278 = {1{`RANDOM}};
  _T_5343_re = _RAND_10278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10279 = {1{`RANDOM}};
  _T_5343_im = _RAND_10279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10280 = {1{`RANDOM}};
  _T_5344_re = _RAND_10280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10281 = {1{`RANDOM}};
  _T_5344_im = _RAND_10281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10282 = {1{`RANDOM}};
  _T_5345_re = _RAND_10282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10283 = {1{`RANDOM}};
  _T_5345_im = _RAND_10283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10284 = {1{`RANDOM}};
  _T_5346_re = _RAND_10284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10285 = {1{`RANDOM}};
  _T_5346_im = _RAND_10285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10286 = {1{`RANDOM}};
  _T_5347_re = _RAND_10286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10287 = {1{`RANDOM}};
  _T_5347_im = _RAND_10287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10288 = {1{`RANDOM}};
  _T_5348_re = _RAND_10288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10289 = {1{`RANDOM}};
  _T_5348_im = _RAND_10289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10290 = {1{`RANDOM}};
  _T_5349_re = _RAND_10290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10291 = {1{`RANDOM}};
  _T_5349_im = _RAND_10291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10292 = {1{`RANDOM}};
  _T_5350_re = _RAND_10292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10293 = {1{`RANDOM}};
  _T_5350_im = _RAND_10293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10294 = {1{`RANDOM}};
  _T_5351_re = _RAND_10294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10295 = {1{`RANDOM}};
  _T_5351_im = _RAND_10295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10296 = {1{`RANDOM}};
  _T_5352_re = _RAND_10296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10297 = {1{`RANDOM}};
  _T_5352_im = _RAND_10297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10298 = {1{`RANDOM}};
  _T_5353_re = _RAND_10298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10299 = {1{`RANDOM}};
  _T_5353_im = _RAND_10299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10300 = {1{`RANDOM}};
  _T_5354_re = _RAND_10300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10301 = {1{`RANDOM}};
  _T_5354_im = _RAND_10301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10302 = {1{`RANDOM}};
  _T_5355_re = _RAND_10302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10303 = {1{`RANDOM}};
  _T_5355_im = _RAND_10303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10304 = {1{`RANDOM}};
  _T_5356_re = _RAND_10304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10305 = {1{`RANDOM}};
  _T_5356_im = _RAND_10305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10306 = {1{`RANDOM}};
  _T_5357_re = _RAND_10306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10307 = {1{`RANDOM}};
  _T_5357_im = _RAND_10307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10308 = {1{`RANDOM}};
  _T_5358_re = _RAND_10308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10309 = {1{`RANDOM}};
  _T_5358_im = _RAND_10309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10310 = {1{`RANDOM}};
  _T_5359_re = _RAND_10310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10311 = {1{`RANDOM}};
  _T_5359_im = _RAND_10311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10312 = {1{`RANDOM}};
  _T_5360_re = _RAND_10312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10313 = {1{`RANDOM}};
  _T_5360_im = _RAND_10313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10314 = {1{`RANDOM}};
  _T_5361_re = _RAND_10314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10315 = {1{`RANDOM}};
  _T_5361_im = _RAND_10315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10316 = {1{`RANDOM}};
  _T_5362_re = _RAND_10316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10317 = {1{`RANDOM}};
  _T_5362_im = _RAND_10317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10318 = {1{`RANDOM}};
  _T_5363_re = _RAND_10318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10319 = {1{`RANDOM}};
  _T_5363_im = _RAND_10319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10320 = {1{`RANDOM}};
  _T_5364_re = _RAND_10320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10321 = {1{`RANDOM}};
  _T_5364_im = _RAND_10321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10322 = {1{`RANDOM}};
  _T_5365_re = _RAND_10322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10323 = {1{`RANDOM}};
  _T_5365_im = _RAND_10323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10324 = {1{`RANDOM}};
  _T_5366_re = _RAND_10324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10325 = {1{`RANDOM}};
  _T_5366_im = _RAND_10325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10326 = {1{`RANDOM}};
  _T_5367_re = _RAND_10326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10327 = {1{`RANDOM}};
  _T_5367_im = _RAND_10327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10328 = {1{`RANDOM}};
  _T_5368_re = _RAND_10328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10329 = {1{`RANDOM}};
  _T_5368_im = _RAND_10329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10330 = {1{`RANDOM}};
  _T_5369_re = _RAND_10330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10331 = {1{`RANDOM}};
  _T_5369_im = _RAND_10331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10332 = {1{`RANDOM}};
  _T_5370_re = _RAND_10332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10333 = {1{`RANDOM}};
  _T_5370_im = _RAND_10333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10334 = {1{`RANDOM}};
  _T_5371_re = _RAND_10334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10335 = {1{`RANDOM}};
  _T_5371_im = _RAND_10335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10336 = {1{`RANDOM}};
  _T_5372_re = _RAND_10336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10337 = {1{`RANDOM}};
  _T_5372_im = _RAND_10337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10338 = {1{`RANDOM}};
  _T_5373_re = _RAND_10338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10339 = {1{`RANDOM}};
  _T_5373_im = _RAND_10339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10340 = {1{`RANDOM}};
  _T_5374_re = _RAND_10340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10341 = {1{`RANDOM}};
  _T_5374_im = _RAND_10341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10342 = {1{`RANDOM}};
  _T_5375_re = _RAND_10342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10343 = {1{`RANDOM}};
  _T_5375_im = _RAND_10343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10344 = {1{`RANDOM}};
  _T_5376_re = _RAND_10344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10345 = {1{`RANDOM}};
  _T_5376_im = _RAND_10345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10346 = {1{`RANDOM}};
  _T_5377_re = _RAND_10346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10347 = {1{`RANDOM}};
  _T_5377_im = _RAND_10347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10348 = {1{`RANDOM}};
  _T_5378_re = _RAND_10348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10349 = {1{`RANDOM}};
  _T_5378_im = _RAND_10349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10350 = {1{`RANDOM}};
  _T_5379_re = _RAND_10350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10351 = {1{`RANDOM}};
  _T_5379_im = _RAND_10351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10352 = {1{`RANDOM}};
  _T_5380_re = _RAND_10352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10353 = {1{`RANDOM}};
  _T_5380_im = _RAND_10353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10354 = {1{`RANDOM}};
  _T_5381_re = _RAND_10354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10355 = {1{`RANDOM}};
  _T_5381_im = _RAND_10355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10356 = {1{`RANDOM}};
  _T_5382_re = _RAND_10356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10357 = {1{`RANDOM}};
  _T_5382_im = _RAND_10357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10358 = {1{`RANDOM}};
  _T_5383_re = _RAND_10358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10359 = {1{`RANDOM}};
  _T_5383_im = _RAND_10359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10360 = {1{`RANDOM}};
  _T_5384_re = _RAND_10360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10361 = {1{`RANDOM}};
  _T_5384_im = _RAND_10361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10362 = {1{`RANDOM}};
  _T_5385_re = _RAND_10362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10363 = {1{`RANDOM}};
  _T_5385_im = _RAND_10363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10364 = {1{`RANDOM}};
  _T_5386_re = _RAND_10364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10365 = {1{`RANDOM}};
  _T_5386_im = _RAND_10365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10366 = {1{`RANDOM}};
  _T_5387_re = _RAND_10366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10367 = {1{`RANDOM}};
  _T_5387_im = _RAND_10367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10368 = {1{`RANDOM}};
  _T_5388_re = _RAND_10368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10369 = {1{`RANDOM}};
  _T_5388_im = _RAND_10369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10370 = {1{`RANDOM}};
  _T_5389_re = _RAND_10370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10371 = {1{`RANDOM}};
  _T_5389_im = _RAND_10371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10372 = {1{`RANDOM}};
  _T_5390_re = _RAND_10372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10373 = {1{`RANDOM}};
  _T_5390_im = _RAND_10373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10374 = {1{`RANDOM}};
  _T_5391_re = _RAND_10374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10375 = {1{`RANDOM}};
  _T_5391_im = _RAND_10375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10376 = {1{`RANDOM}};
  _T_5392_re = _RAND_10376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10377 = {1{`RANDOM}};
  _T_5392_im = _RAND_10377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10378 = {1{`RANDOM}};
  _T_5393_re = _RAND_10378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10379 = {1{`RANDOM}};
  _T_5393_im = _RAND_10379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10380 = {1{`RANDOM}};
  _T_5394_re = _RAND_10380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10381 = {1{`RANDOM}};
  _T_5394_im = _RAND_10381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10382 = {1{`RANDOM}};
  _T_5395_re = _RAND_10382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10383 = {1{`RANDOM}};
  _T_5395_im = _RAND_10383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10384 = {1{`RANDOM}};
  _T_5396_re = _RAND_10384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10385 = {1{`RANDOM}};
  _T_5396_im = _RAND_10385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10386 = {1{`RANDOM}};
  _T_5397_re = _RAND_10386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10387 = {1{`RANDOM}};
  _T_5397_im = _RAND_10387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10388 = {1{`RANDOM}};
  _T_5398_re = _RAND_10388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10389 = {1{`RANDOM}};
  _T_5398_im = _RAND_10389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10390 = {1{`RANDOM}};
  _T_5399_re = _RAND_10390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10391 = {1{`RANDOM}};
  _T_5399_im = _RAND_10391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10392 = {1{`RANDOM}};
  _T_5400_re = _RAND_10392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10393 = {1{`RANDOM}};
  _T_5400_im = _RAND_10393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10394 = {1{`RANDOM}};
  _T_5401_re = _RAND_10394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10395 = {1{`RANDOM}};
  _T_5401_im = _RAND_10395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10396 = {1{`RANDOM}};
  _T_5402_re = _RAND_10396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10397 = {1{`RANDOM}};
  _T_5402_im = _RAND_10397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10398 = {1{`RANDOM}};
  _T_5403_re = _RAND_10398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10399 = {1{`RANDOM}};
  _T_5403_im = _RAND_10399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10400 = {1{`RANDOM}};
  _T_5404_re = _RAND_10400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10401 = {1{`RANDOM}};
  _T_5404_im = _RAND_10401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10402 = {1{`RANDOM}};
  _T_5405_re = _RAND_10402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10403 = {1{`RANDOM}};
  _T_5405_im = _RAND_10403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10404 = {1{`RANDOM}};
  _T_5406_re = _RAND_10404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10405 = {1{`RANDOM}};
  _T_5406_im = _RAND_10405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10406 = {1{`RANDOM}};
  _T_5407_re = _RAND_10406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10407 = {1{`RANDOM}};
  _T_5407_im = _RAND_10407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10408 = {1{`RANDOM}};
  _T_5408_re = _RAND_10408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10409 = {1{`RANDOM}};
  _T_5408_im = _RAND_10409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10410 = {1{`RANDOM}};
  _T_5409_re = _RAND_10410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10411 = {1{`RANDOM}};
  _T_5409_im = _RAND_10411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10412 = {1{`RANDOM}};
  _T_5410_re = _RAND_10412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10413 = {1{`RANDOM}};
  _T_5410_im = _RAND_10413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10414 = {1{`RANDOM}};
  _T_5411_re = _RAND_10414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10415 = {1{`RANDOM}};
  _T_5411_im = _RAND_10415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10416 = {1{`RANDOM}};
  _T_5412_re = _RAND_10416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10417 = {1{`RANDOM}};
  _T_5412_im = _RAND_10417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10418 = {1{`RANDOM}};
  _T_5413_re = _RAND_10418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10419 = {1{`RANDOM}};
  _T_5413_im = _RAND_10419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10420 = {1{`RANDOM}};
  _T_5414_re = _RAND_10420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10421 = {1{`RANDOM}};
  _T_5414_im = _RAND_10421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10422 = {1{`RANDOM}};
  _T_5415_re = _RAND_10422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10423 = {1{`RANDOM}};
  _T_5415_im = _RAND_10423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10424 = {1{`RANDOM}};
  _T_5416_re = _RAND_10424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10425 = {1{`RANDOM}};
  _T_5416_im = _RAND_10425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10426 = {1{`RANDOM}};
  _T_5417_re = _RAND_10426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10427 = {1{`RANDOM}};
  _T_5417_im = _RAND_10427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10428 = {1{`RANDOM}};
  _T_5418_re = _RAND_10428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10429 = {1{`RANDOM}};
  _T_5418_im = _RAND_10429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10430 = {1{`RANDOM}};
  _T_5419_re = _RAND_10430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10431 = {1{`RANDOM}};
  _T_5419_im = _RAND_10431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10432 = {1{`RANDOM}};
  _T_5420_re = _RAND_10432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10433 = {1{`RANDOM}};
  _T_5420_im = _RAND_10433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10434 = {1{`RANDOM}};
  _T_5421_re = _RAND_10434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10435 = {1{`RANDOM}};
  _T_5421_im = _RAND_10435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10436 = {1{`RANDOM}};
  _T_5422_re = _RAND_10436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10437 = {1{`RANDOM}};
  _T_5422_im = _RAND_10437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10438 = {1{`RANDOM}};
  _T_5423_re = _RAND_10438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10439 = {1{`RANDOM}};
  _T_5423_im = _RAND_10439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10440 = {1{`RANDOM}};
  _T_5424_re = _RAND_10440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10441 = {1{`RANDOM}};
  _T_5424_im = _RAND_10441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10442 = {1{`RANDOM}};
  _T_5425_re = _RAND_10442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10443 = {1{`RANDOM}};
  _T_5425_im = _RAND_10443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10444 = {1{`RANDOM}};
  _T_5426_re = _RAND_10444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10445 = {1{`RANDOM}};
  _T_5426_im = _RAND_10445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10446 = {1{`RANDOM}};
  _T_5427_re = _RAND_10446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10447 = {1{`RANDOM}};
  _T_5427_im = _RAND_10447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10448 = {1{`RANDOM}};
  _T_5428_re = _RAND_10448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10449 = {1{`RANDOM}};
  _T_5428_im = _RAND_10449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10450 = {1{`RANDOM}};
  _T_5429_re = _RAND_10450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10451 = {1{`RANDOM}};
  _T_5429_im = _RAND_10451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10452 = {1{`RANDOM}};
  _T_5430_re = _RAND_10452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10453 = {1{`RANDOM}};
  _T_5430_im = _RAND_10453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10454 = {1{`RANDOM}};
  _T_5431_re = _RAND_10454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10455 = {1{`RANDOM}};
  _T_5431_im = _RAND_10455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10456 = {1{`RANDOM}};
  _T_5432_re = _RAND_10456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10457 = {1{`RANDOM}};
  _T_5432_im = _RAND_10457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10458 = {1{`RANDOM}};
  _T_5433_re = _RAND_10458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10459 = {1{`RANDOM}};
  _T_5433_im = _RAND_10459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10460 = {1{`RANDOM}};
  _T_5434_re = _RAND_10460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10461 = {1{`RANDOM}};
  _T_5434_im = _RAND_10461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10462 = {1{`RANDOM}};
  _T_5435_re = _RAND_10462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10463 = {1{`RANDOM}};
  _T_5435_im = _RAND_10463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10464 = {1{`RANDOM}};
  _T_5436_re = _RAND_10464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10465 = {1{`RANDOM}};
  _T_5436_im = _RAND_10465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10466 = {1{`RANDOM}};
  _T_5437_re = _RAND_10466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10467 = {1{`RANDOM}};
  _T_5437_im = _RAND_10467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10468 = {1{`RANDOM}};
  _T_5438_re = _RAND_10468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10469 = {1{`RANDOM}};
  _T_5438_im = _RAND_10469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10470 = {1{`RANDOM}};
  _T_5439_re = _RAND_10470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10471 = {1{`RANDOM}};
  _T_5439_im = _RAND_10471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10472 = {1{`RANDOM}};
  _T_5440_re = _RAND_10472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10473 = {1{`RANDOM}};
  _T_5440_im = _RAND_10473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10474 = {1{`RANDOM}};
  _T_5441_re = _RAND_10474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10475 = {1{`RANDOM}};
  _T_5441_im = _RAND_10475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10476 = {1{`RANDOM}};
  _T_5442_re = _RAND_10476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10477 = {1{`RANDOM}};
  _T_5442_im = _RAND_10477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10478 = {1{`RANDOM}};
  _T_5443_re = _RAND_10478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10479 = {1{`RANDOM}};
  _T_5443_im = _RAND_10479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10480 = {1{`RANDOM}};
  _T_5444_re = _RAND_10480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10481 = {1{`RANDOM}};
  _T_5444_im = _RAND_10481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10482 = {1{`RANDOM}};
  _T_5445_re = _RAND_10482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10483 = {1{`RANDOM}};
  _T_5445_im = _RAND_10483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10484 = {1{`RANDOM}};
  _T_5446_re = _RAND_10484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10485 = {1{`RANDOM}};
  _T_5446_im = _RAND_10485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10486 = {1{`RANDOM}};
  _T_5447_re = _RAND_10486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10487 = {1{`RANDOM}};
  _T_5447_im = _RAND_10487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10488 = {1{`RANDOM}};
  _T_5448_re = _RAND_10488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10489 = {1{`RANDOM}};
  _T_5448_im = _RAND_10489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10490 = {1{`RANDOM}};
  _T_5449_re = _RAND_10490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10491 = {1{`RANDOM}};
  _T_5449_im = _RAND_10491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10492 = {1{`RANDOM}};
  _T_5450_re = _RAND_10492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10493 = {1{`RANDOM}};
  _T_5450_im = _RAND_10493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10494 = {1{`RANDOM}};
  _T_5451_re = _RAND_10494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10495 = {1{`RANDOM}};
  _T_5451_im = _RAND_10495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10496 = {1{`RANDOM}};
  _T_5452_re = _RAND_10496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10497 = {1{`RANDOM}};
  _T_5452_im = _RAND_10497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10498 = {1{`RANDOM}};
  _T_5453_re = _RAND_10498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10499 = {1{`RANDOM}};
  _T_5453_im = _RAND_10499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10500 = {1{`RANDOM}};
  _T_5454_re = _RAND_10500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10501 = {1{`RANDOM}};
  _T_5454_im = _RAND_10501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10502 = {1{`RANDOM}};
  _T_5455_re = _RAND_10502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10503 = {1{`RANDOM}};
  _T_5455_im = _RAND_10503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10504 = {1{`RANDOM}};
  _T_5456_re = _RAND_10504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10505 = {1{`RANDOM}};
  _T_5456_im = _RAND_10505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10506 = {1{`RANDOM}};
  _T_5457_re = _RAND_10506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10507 = {1{`RANDOM}};
  _T_5457_im = _RAND_10507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10508 = {1{`RANDOM}};
  _T_5458_re = _RAND_10508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10509 = {1{`RANDOM}};
  _T_5458_im = _RAND_10509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10510 = {1{`RANDOM}};
  _T_5459_re = _RAND_10510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10511 = {1{`RANDOM}};
  _T_5459_im = _RAND_10511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10512 = {1{`RANDOM}};
  _T_5460_re = _RAND_10512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10513 = {1{`RANDOM}};
  _T_5460_im = _RAND_10513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10514 = {1{`RANDOM}};
  _T_5461_re = _RAND_10514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10515 = {1{`RANDOM}};
  _T_5461_im = _RAND_10515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10516 = {1{`RANDOM}};
  _T_5462_re = _RAND_10516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10517 = {1{`RANDOM}};
  _T_5462_im = _RAND_10517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10518 = {1{`RANDOM}};
  _T_5463_re = _RAND_10518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10519 = {1{`RANDOM}};
  _T_5463_im = _RAND_10519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10520 = {1{`RANDOM}};
  _T_5464_re = _RAND_10520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10521 = {1{`RANDOM}};
  _T_5464_im = _RAND_10521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10522 = {1{`RANDOM}};
  _T_5465_re = _RAND_10522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10523 = {1{`RANDOM}};
  _T_5465_im = _RAND_10523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10524 = {1{`RANDOM}};
  _T_5466_re = _RAND_10524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10525 = {1{`RANDOM}};
  _T_5466_im = _RAND_10525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10526 = {1{`RANDOM}};
  _T_5467_re = _RAND_10526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10527 = {1{`RANDOM}};
  _T_5467_im = _RAND_10527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10528 = {1{`RANDOM}};
  _T_5468_re = _RAND_10528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10529 = {1{`RANDOM}};
  _T_5468_im = _RAND_10529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10530 = {1{`RANDOM}};
  _T_5469_re = _RAND_10530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10531 = {1{`RANDOM}};
  _T_5469_im = _RAND_10531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10532 = {1{`RANDOM}};
  _T_5470_re = _RAND_10532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10533 = {1{`RANDOM}};
  _T_5470_im = _RAND_10533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10534 = {1{`RANDOM}};
  _T_5471_re = _RAND_10534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10535 = {1{`RANDOM}};
  _T_5471_im = _RAND_10535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10536 = {1{`RANDOM}};
  _T_5472_re = _RAND_10536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10537 = {1{`RANDOM}};
  _T_5472_im = _RAND_10537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10538 = {1{`RANDOM}};
  _T_5473_re = _RAND_10538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10539 = {1{`RANDOM}};
  _T_5473_im = _RAND_10539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10540 = {1{`RANDOM}};
  _T_5474_re = _RAND_10540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10541 = {1{`RANDOM}};
  _T_5474_im = _RAND_10541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10542 = {1{`RANDOM}};
  _T_5475_re = _RAND_10542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10543 = {1{`RANDOM}};
  _T_5475_im = _RAND_10543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10544 = {1{`RANDOM}};
  _T_5476_re = _RAND_10544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10545 = {1{`RANDOM}};
  _T_5476_im = _RAND_10545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10546 = {1{`RANDOM}};
  _T_5477_re = _RAND_10546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10547 = {1{`RANDOM}};
  _T_5477_im = _RAND_10547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10548 = {1{`RANDOM}};
  _T_5478_re = _RAND_10548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10549 = {1{`RANDOM}};
  _T_5478_im = _RAND_10549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10550 = {1{`RANDOM}};
  _T_5479_re = _RAND_10550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10551 = {1{`RANDOM}};
  _T_5479_im = _RAND_10551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10552 = {1{`RANDOM}};
  _T_5480_re = _RAND_10552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10553 = {1{`RANDOM}};
  _T_5480_im = _RAND_10553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10554 = {1{`RANDOM}};
  _T_5481_re = _RAND_10554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10555 = {1{`RANDOM}};
  _T_5481_im = _RAND_10555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10556 = {1{`RANDOM}};
  _T_5482_re = _RAND_10556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10557 = {1{`RANDOM}};
  _T_5482_im = _RAND_10557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10558 = {1{`RANDOM}};
  _T_5483_re = _RAND_10558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10559 = {1{`RANDOM}};
  _T_5483_im = _RAND_10559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10560 = {1{`RANDOM}};
  _T_5484_re = _RAND_10560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10561 = {1{`RANDOM}};
  _T_5484_im = _RAND_10561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10562 = {1{`RANDOM}};
  _T_5485_re = _RAND_10562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10563 = {1{`RANDOM}};
  _T_5485_im = _RAND_10563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10564 = {1{`RANDOM}};
  _T_5486_re = _RAND_10564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10565 = {1{`RANDOM}};
  _T_5486_im = _RAND_10565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10566 = {1{`RANDOM}};
  _T_5487_re = _RAND_10566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10567 = {1{`RANDOM}};
  _T_5487_im = _RAND_10567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10568 = {1{`RANDOM}};
  _T_5488_re = _RAND_10568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10569 = {1{`RANDOM}};
  _T_5488_im = _RAND_10569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10570 = {1{`RANDOM}};
  _T_5489_re = _RAND_10570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10571 = {1{`RANDOM}};
  _T_5489_im = _RAND_10571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10572 = {1{`RANDOM}};
  _T_5490_re = _RAND_10572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10573 = {1{`RANDOM}};
  _T_5490_im = _RAND_10573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10574 = {1{`RANDOM}};
  _T_5491_re = _RAND_10574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10575 = {1{`RANDOM}};
  _T_5491_im = _RAND_10575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10576 = {1{`RANDOM}};
  _T_5492_re = _RAND_10576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10577 = {1{`RANDOM}};
  _T_5492_im = _RAND_10577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10578 = {1{`RANDOM}};
  _T_5493_re = _RAND_10578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10579 = {1{`RANDOM}};
  _T_5493_im = _RAND_10579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10580 = {1{`RANDOM}};
  _T_5494_re = _RAND_10580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10581 = {1{`RANDOM}};
  _T_5494_im = _RAND_10581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10582 = {1{`RANDOM}};
  _T_5495_re = _RAND_10582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10583 = {1{`RANDOM}};
  _T_5495_im = _RAND_10583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10584 = {1{`RANDOM}};
  _T_5496_re = _RAND_10584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10585 = {1{`RANDOM}};
  _T_5496_im = _RAND_10585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10586 = {1{`RANDOM}};
  _T_5497_re = _RAND_10586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10587 = {1{`RANDOM}};
  _T_5497_im = _RAND_10587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10588 = {1{`RANDOM}};
  _T_5498_re = _RAND_10588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10589 = {1{`RANDOM}};
  _T_5498_im = _RAND_10589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10590 = {1{`RANDOM}};
  _T_5499_re = _RAND_10590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10591 = {1{`RANDOM}};
  _T_5499_im = _RAND_10591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10592 = {1{`RANDOM}};
  _T_5500_re = _RAND_10592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10593 = {1{`RANDOM}};
  _T_5500_im = _RAND_10593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10594 = {1{`RANDOM}};
  _T_5501_re = _RAND_10594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10595 = {1{`RANDOM}};
  _T_5501_im = _RAND_10595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10596 = {1{`RANDOM}};
  _T_5502_re = _RAND_10596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10597 = {1{`RANDOM}};
  _T_5502_im = _RAND_10597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10598 = {1{`RANDOM}};
  _T_5503_re = _RAND_10598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10599 = {1{`RANDOM}};
  _T_5503_im = _RAND_10599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10600 = {1{`RANDOM}};
  _T_5504_re = _RAND_10600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10601 = {1{`RANDOM}};
  _T_5504_im = _RAND_10601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10602 = {1{`RANDOM}};
  _T_5505_re = _RAND_10602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10603 = {1{`RANDOM}};
  _T_5505_im = _RAND_10603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10604 = {1{`RANDOM}};
  _T_5506_re = _RAND_10604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10605 = {1{`RANDOM}};
  _T_5506_im = _RAND_10605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10606 = {1{`RANDOM}};
  _T_5507_re = _RAND_10606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10607 = {1{`RANDOM}};
  _T_5507_im = _RAND_10607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10608 = {1{`RANDOM}};
  _T_5508_re = _RAND_10608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10609 = {1{`RANDOM}};
  _T_5508_im = _RAND_10609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10610 = {1{`RANDOM}};
  _T_5509_re = _RAND_10610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10611 = {1{`RANDOM}};
  _T_5509_im = _RAND_10611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10612 = {1{`RANDOM}};
  _T_5510_re = _RAND_10612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10613 = {1{`RANDOM}};
  _T_5510_im = _RAND_10613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10614 = {1{`RANDOM}};
  _T_5511_re = _RAND_10614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10615 = {1{`RANDOM}};
  _T_5511_im = _RAND_10615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10616 = {1{`RANDOM}};
  _T_5512_re = _RAND_10616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10617 = {1{`RANDOM}};
  _T_5512_im = _RAND_10617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10618 = {1{`RANDOM}};
  _T_5513_re = _RAND_10618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10619 = {1{`RANDOM}};
  _T_5513_im = _RAND_10619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10620 = {1{`RANDOM}};
  _T_5514_re = _RAND_10620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10621 = {1{`RANDOM}};
  _T_5514_im = _RAND_10621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10622 = {1{`RANDOM}};
  _T_5515_re = _RAND_10622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10623 = {1{`RANDOM}};
  _T_5515_im = _RAND_10623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10624 = {1{`RANDOM}};
  _T_5516_re = _RAND_10624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10625 = {1{`RANDOM}};
  _T_5516_im = _RAND_10625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10626 = {1{`RANDOM}};
  _T_5517_re = _RAND_10626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10627 = {1{`RANDOM}};
  _T_5517_im = _RAND_10627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10628 = {1{`RANDOM}};
  _T_5518_re = _RAND_10628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10629 = {1{`RANDOM}};
  _T_5518_im = _RAND_10629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10630 = {1{`RANDOM}};
  _T_5519_re = _RAND_10630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10631 = {1{`RANDOM}};
  _T_5519_im = _RAND_10631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10632 = {1{`RANDOM}};
  _T_5520_re = _RAND_10632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10633 = {1{`RANDOM}};
  _T_5520_im = _RAND_10633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10634 = {1{`RANDOM}};
  _T_5521_re = _RAND_10634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10635 = {1{`RANDOM}};
  _T_5521_im = _RAND_10635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10636 = {1{`RANDOM}};
  _T_5522_re = _RAND_10636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10637 = {1{`RANDOM}};
  _T_5522_im = _RAND_10637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10638 = {1{`RANDOM}};
  _T_5523_re = _RAND_10638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10639 = {1{`RANDOM}};
  _T_5523_im = _RAND_10639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10640 = {1{`RANDOM}};
  _T_5524_re = _RAND_10640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10641 = {1{`RANDOM}};
  _T_5524_im = _RAND_10641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10642 = {1{`RANDOM}};
  _T_5525_re = _RAND_10642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10643 = {1{`RANDOM}};
  _T_5525_im = _RAND_10643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10644 = {1{`RANDOM}};
  _T_5526_re = _RAND_10644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10645 = {1{`RANDOM}};
  _T_5526_im = _RAND_10645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10646 = {1{`RANDOM}};
  _T_5527_re = _RAND_10646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10647 = {1{`RANDOM}};
  _T_5527_im = _RAND_10647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10648 = {1{`RANDOM}};
  _T_5528_re = _RAND_10648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10649 = {1{`RANDOM}};
  _T_5528_im = _RAND_10649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10650 = {1{`RANDOM}};
  _T_5529_re = _RAND_10650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10651 = {1{`RANDOM}};
  _T_5529_im = _RAND_10651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10652 = {1{`RANDOM}};
  _T_5530_re = _RAND_10652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10653 = {1{`RANDOM}};
  _T_5530_im = _RAND_10653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10654 = {1{`RANDOM}};
  _T_5531_re = _RAND_10654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10655 = {1{`RANDOM}};
  _T_5531_im = _RAND_10655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10656 = {1{`RANDOM}};
  _T_5532_re = _RAND_10656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10657 = {1{`RANDOM}};
  _T_5532_im = _RAND_10657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10658 = {1{`RANDOM}};
  _T_5533_re = _RAND_10658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10659 = {1{`RANDOM}};
  _T_5533_im = _RAND_10659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10660 = {1{`RANDOM}};
  _T_5534_re = _RAND_10660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10661 = {1{`RANDOM}};
  _T_5534_im = _RAND_10661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10662 = {1{`RANDOM}};
  _T_5535_re = _RAND_10662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10663 = {1{`RANDOM}};
  _T_5535_im = _RAND_10663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10664 = {1{`RANDOM}};
  _T_5536_re = _RAND_10664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10665 = {1{`RANDOM}};
  _T_5536_im = _RAND_10665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10666 = {1{`RANDOM}};
  _T_5537_re = _RAND_10666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10667 = {1{`RANDOM}};
  _T_5537_im = _RAND_10667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10668 = {1{`RANDOM}};
  _T_5538_re = _RAND_10668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10669 = {1{`RANDOM}};
  _T_5538_im = _RAND_10669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10670 = {1{`RANDOM}};
  _T_5539_re = _RAND_10670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10671 = {1{`RANDOM}};
  _T_5539_im = _RAND_10671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10672 = {1{`RANDOM}};
  _T_5540_re = _RAND_10672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10673 = {1{`RANDOM}};
  _T_5540_im = _RAND_10673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10674 = {1{`RANDOM}};
  _T_5541_re = _RAND_10674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10675 = {1{`RANDOM}};
  _T_5541_im = _RAND_10675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10676 = {1{`RANDOM}};
  _T_5542_re = _RAND_10676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10677 = {1{`RANDOM}};
  _T_5542_im = _RAND_10677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10678 = {1{`RANDOM}};
  _T_5543_re = _RAND_10678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10679 = {1{`RANDOM}};
  _T_5543_im = _RAND_10679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10680 = {1{`RANDOM}};
  _T_5544_re = _RAND_10680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10681 = {1{`RANDOM}};
  _T_5544_im = _RAND_10681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10682 = {1{`RANDOM}};
  _T_5545_re = _RAND_10682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10683 = {1{`RANDOM}};
  _T_5545_im = _RAND_10683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10684 = {1{`RANDOM}};
  _T_5546_re = _RAND_10684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10685 = {1{`RANDOM}};
  _T_5546_im = _RAND_10685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10686 = {1{`RANDOM}};
  _T_5547_re = _RAND_10686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10687 = {1{`RANDOM}};
  _T_5547_im = _RAND_10687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10688 = {1{`RANDOM}};
  _T_5548_re = _RAND_10688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10689 = {1{`RANDOM}};
  _T_5548_im = _RAND_10689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10690 = {1{`RANDOM}};
  _T_5549_re = _RAND_10690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10691 = {1{`RANDOM}};
  _T_5549_im = _RAND_10691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10692 = {1{`RANDOM}};
  _T_5550_re = _RAND_10692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10693 = {1{`RANDOM}};
  _T_5550_im = _RAND_10693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10694 = {1{`RANDOM}};
  _T_5551_re = _RAND_10694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10695 = {1{`RANDOM}};
  _T_5551_im = _RAND_10695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10696 = {1{`RANDOM}};
  _T_5552_re = _RAND_10696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10697 = {1{`RANDOM}};
  _T_5552_im = _RAND_10697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10698 = {1{`RANDOM}};
  _T_5553_re = _RAND_10698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10699 = {1{`RANDOM}};
  _T_5553_im = _RAND_10699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10700 = {1{`RANDOM}};
  _T_5554_re = _RAND_10700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10701 = {1{`RANDOM}};
  _T_5554_im = _RAND_10701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10702 = {1{`RANDOM}};
  _T_5555_re = _RAND_10702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10703 = {1{`RANDOM}};
  _T_5555_im = _RAND_10703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10704 = {1{`RANDOM}};
  _T_5556_re = _RAND_10704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10705 = {1{`RANDOM}};
  _T_5556_im = _RAND_10705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10706 = {1{`RANDOM}};
  _T_5557_re = _RAND_10706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10707 = {1{`RANDOM}};
  _T_5557_im = _RAND_10707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10708 = {1{`RANDOM}};
  _T_5558_re = _RAND_10708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10709 = {1{`RANDOM}};
  _T_5558_im = _RAND_10709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10710 = {1{`RANDOM}};
  _T_5559_re = _RAND_10710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10711 = {1{`RANDOM}};
  _T_5559_im = _RAND_10711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10712 = {1{`RANDOM}};
  _T_5560_re = _RAND_10712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10713 = {1{`RANDOM}};
  _T_5560_im = _RAND_10713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10714 = {1{`RANDOM}};
  _T_5561_re = _RAND_10714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10715 = {1{`RANDOM}};
  _T_5561_im = _RAND_10715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10716 = {1{`RANDOM}};
  _T_5562_re = _RAND_10716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10717 = {1{`RANDOM}};
  _T_5562_im = _RAND_10717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10718 = {1{`RANDOM}};
  _T_5563_re = _RAND_10718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10719 = {1{`RANDOM}};
  _T_5563_im = _RAND_10719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10720 = {1{`RANDOM}};
  _T_5564_re = _RAND_10720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10721 = {1{`RANDOM}};
  _T_5564_im = _RAND_10721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10722 = {1{`RANDOM}};
  _T_5565_re = _RAND_10722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10723 = {1{`RANDOM}};
  _T_5565_im = _RAND_10723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10724 = {1{`RANDOM}};
  _T_5566_re = _RAND_10724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10725 = {1{`RANDOM}};
  _T_5566_im = _RAND_10725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10726 = {1{`RANDOM}};
  _T_5567_re = _RAND_10726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10727 = {1{`RANDOM}};
  _T_5567_im = _RAND_10727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10728 = {1{`RANDOM}};
  _T_5568_re = _RAND_10728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10729 = {1{`RANDOM}};
  _T_5568_im = _RAND_10729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10730 = {1{`RANDOM}};
  _T_5569_re = _RAND_10730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10731 = {1{`RANDOM}};
  _T_5569_im = _RAND_10731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10732 = {1{`RANDOM}};
  _T_5570_re = _RAND_10732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10733 = {1{`RANDOM}};
  _T_5570_im = _RAND_10733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10734 = {1{`RANDOM}};
  _T_5571_re = _RAND_10734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10735 = {1{`RANDOM}};
  _T_5571_im = _RAND_10735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10736 = {1{`RANDOM}};
  _T_5572_re = _RAND_10736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10737 = {1{`RANDOM}};
  _T_5572_im = _RAND_10737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10738 = {1{`RANDOM}};
  _T_5573_re = _RAND_10738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10739 = {1{`RANDOM}};
  _T_5573_im = _RAND_10739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10740 = {1{`RANDOM}};
  _T_5574_re = _RAND_10740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10741 = {1{`RANDOM}};
  _T_5574_im = _RAND_10741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10742 = {1{`RANDOM}};
  _T_5575_re = _RAND_10742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10743 = {1{`RANDOM}};
  _T_5575_im = _RAND_10743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10744 = {1{`RANDOM}};
  _T_5576_re = _RAND_10744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10745 = {1{`RANDOM}};
  _T_5576_im = _RAND_10745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10746 = {1{`RANDOM}};
  _T_5577_re = _RAND_10746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10747 = {1{`RANDOM}};
  _T_5577_im = _RAND_10747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10748 = {1{`RANDOM}};
  _T_5578_re = _RAND_10748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10749 = {1{`RANDOM}};
  _T_5578_im = _RAND_10749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10750 = {1{`RANDOM}};
  _T_5579_re = _RAND_10750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10751 = {1{`RANDOM}};
  _T_5579_im = _RAND_10751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10752 = {1{`RANDOM}};
  _T_5580_re = _RAND_10752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10753 = {1{`RANDOM}};
  _T_5580_im = _RAND_10753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10754 = {1{`RANDOM}};
  _T_5586_re = _RAND_10754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10755 = {1{`RANDOM}};
  _T_5586_im = _RAND_10755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10756 = {1{`RANDOM}};
  _T_5587_re = _RAND_10756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10757 = {1{`RANDOM}};
  _T_5587_im = _RAND_10757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10758 = {1{`RANDOM}};
  _T_5588_re = _RAND_10758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10759 = {1{`RANDOM}};
  _T_5588_im = _RAND_10759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10760 = {1{`RANDOM}};
  _T_5589_re = _RAND_10760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10761 = {1{`RANDOM}};
  _T_5589_im = _RAND_10761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10762 = {1{`RANDOM}};
  _T_5590_re = _RAND_10762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10763 = {1{`RANDOM}};
  _T_5590_im = _RAND_10763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10764 = {1{`RANDOM}};
  _T_5591_re = _RAND_10764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10765 = {1{`RANDOM}};
  _T_5591_im = _RAND_10765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10766 = {1{`RANDOM}};
  _T_5592_re = _RAND_10766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10767 = {1{`RANDOM}};
  _T_5592_im = _RAND_10767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10768 = {1{`RANDOM}};
  _T_5593_re = _RAND_10768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10769 = {1{`RANDOM}};
  _T_5593_im = _RAND_10769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10770 = {1{`RANDOM}};
  _T_5594_re = _RAND_10770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10771 = {1{`RANDOM}};
  _T_5594_im = _RAND_10771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10772 = {1{`RANDOM}};
  _T_5595_re = _RAND_10772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10773 = {1{`RANDOM}};
  _T_5595_im = _RAND_10773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10774 = {1{`RANDOM}};
  _T_5596_re = _RAND_10774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10775 = {1{`RANDOM}};
  _T_5596_im = _RAND_10775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10776 = {1{`RANDOM}};
  _T_5597_re = _RAND_10776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10777 = {1{`RANDOM}};
  _T_5597_im = _RAND_10777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10778 = {1{`RANDOM}};
  _T_5598_re = _RAND_10778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10779 = {1{`RANDOM}};
  _T_5598_im = _RAND_10779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10780 = {1{`RANDOM}};
  _T_5599_re = _RAND_10780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10781 = {1{`RANDOM}};
  _T_5599_im = _RAND_10781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10782 = {1{`RANDOM}};
  _T_5600_re = _RAND_10782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10783 = {1{`RANDOM}};
  _T_5600_im = _RAND_10783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10784 = {1{`RANDOM}};
  _T_5601_re = _RAND_10784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10785 = {1{`RANDOM}};
  _T_5601_im = _RAND_10785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10786 = {1{`RANDOM}};
  _T_5602_re = _RAND_10786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10787 = {1{`RANDOM}};
  _T_5602_im = _RAND_10787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10788 = {1{`RANDOM}};
  _T_5603_re = _RAND_10788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10789 = {1{`RANDOM}};
  _T_5603_im = _RAND_10789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10790 = {1{`RANDOM}};
  _T_5604_re = _RAND_10790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10791 = {1{`RANDOM}};
  _T_5604_im = _RAND_10791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10792 = {1{`RANDOM}};
  _T_5605_re = _RAND_10792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10793 = {1{`RANDOM}};
  _T_5605_im = _RAND_10793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10794 = {1{`RANDOM}};
  _T_5606_re = _RAND_10794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10795 = {1{`RANDOM}};
  _T_5606_im = _RAND_10795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10796 = {1{`RANDOM}};
  _T_5607_re = _RAND_10796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10797 = {1{`RANDOM}};
  _T_5607_im = _RAND_10797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10798 = {1{`RANDOM}};
  _T_5608_re = _RAND_10798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10799 = {1{`RANDOM}};
  _T_5608_im = _RAND_10799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10800 = {1{`RANDOM}};
  _T_5609_re = _RAND_10800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10801 = {1{`RANDOM}};
  _T_5609_im = _RAND_10801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10802 = {1{`RANDOM}};
  _T_5610_re = _RAND_10802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10803 = {1{`RANDOM}};
  _T_5610_im = _RAND_10803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10804 = {1{`RANDOM}};
  _T_5611_re = _RAND_10804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10805 = {1{`RANDOM}};
  _T_5611_im = _RAND_10805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10806 = {1{`RANDOM}};
  _T_5612_re = _RAND_10806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10807 = {1{`RANDOM}};
  _T_5612_im = _RAND_10807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10808 = {1{`RANDOM}};
  _T_5613_re = _RAND_10808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10809 = {1{`RANDOM}};
  _T_5613_im = _RAND_10809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10810 = {1{`RANDOM}};
  _T_5614_re = _RAND_10810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10811 = {1{`RANDOM}};
  _T_5614_im = _RAND_10811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10812 = {1{`RANDOM}};
  _T_5615_re = _RAND_10812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10813 = {1{`RANDOM}};
  _T_5615_im = _RAND_10813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10814 = {1{`RANDOM}};
  _T_5616_re = _RAND_10814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10815 = {1{`RANDOM}};
  _T_5616_im = _RAND_10815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10816 = {1{`RANDOM}};
  _T_5617_re = _RAND_10816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10817 = {1{`RANDOM}};
  _T_5617_im = _RAND_10817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10818 = {1{`RANDOM}};
  _T_5618_re = _RAND_10818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10819 = {1{`RANDOM}};
  _T_5618_im = _RAND_10819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10820 = {1{`RANDOM}};
  _T_5619_re = _RAND_10820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10821 = {1{`RANDOM}};
  _T_5619_im = _RAND_10821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10822 = {1{`RANDOM}};
  _T_5620_re = _RAND_10822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10823 = {1{`RANDOM}};
  _T_5620_im = _RAND_10823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10824 = {1{`RANDOM}};
  _T_5621_re = _RAND_10824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10825 = {1{`RANDOM}};
  _T_5621_im = _RAND_10825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10826 = {1{`RANDOM}};
  _T_5622_re = _RAND_10826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10827 = {1{`RANDOM}};
  _T_5622_im = _RAND_10827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10828 = {1{`RANDOM}};
  _T_5623_re = _RAND_10828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10829 = {1{`RANDOM}};
  _T_5623_im = _RAND_10829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10830 = {1{`RANDOM}};
  _T_5624_re = _RAND_10830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10831 = {1{`RANDOM}};
  _T_5624_im = _RAND_10831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10832 = {1{`RANDOM}};
  _T_5625_re = _RAND_10832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10833 = {1{`RANDOM}};
  _T_5625_im = _RAND_10833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10834 = {1{`RANDOM}};
  _T_5626_re = _RAND_10834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10835 = {1{`RANDOM}};
  _T_5626_im = _RAND_10835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10836 = {1{`RANDOM}};
  _T_5627_re = _RAND_10836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10837 = {1{`RANDOM}};
  _T_5627_im = _RAND_10837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10838 = {1{`RANDOM}};
  _T_5628_re = _RAND_10838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10839 = {1{`RANDOM}};
  _T_5628_im = _RAND_10839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10840 = {1{`RANDOM}};
  _T_5629_re = _RAND_10840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10841 = {1{`RANDOM}};
  _T_5629_im = _RAND_10841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10842 = {1{`RANDOM}};
  _T_5630_re = _RAND_10842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10843 = {1{`RANDOM}};
  _T_5630_im = _RAND_10843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10844 = {1{`RANDOM}};
  _T_5631_re = _RAND_10844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10845 = {1{`RANDOM}};
  _T_5631_im = _RAND_10845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10846 = {1{`RANDOM}};
  _T_5632_re = _RAND_10846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10847 = {1{`RANDOM}};
  _T_5632_im = _RAND_10847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10848 = {1{`RANDOM}};
  _T_5633_re = _RAND_10848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10849 = {1{`RANDOM}};
  _T_5633_im = _RAND_10849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10850 = {1{`RANDOM}};
  _T_5634_re = _RAND_10850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10851 = {1{`RANDOM}};
  _T_5634_im = _RAND_10851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10852 = {1{`RANDOM}};
  _T_5635_re = _RAND_10852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10853 = {1{`RANDOM}};
  _T_5635_im = _RAND_10853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10854 = {1{`RANDOM}};
  _T_5636_re = _RAND_10854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10855 = {1{`RANDOM}};
  _T_5636_im = _RAND_10855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10856 = {1{`RANDOM}};
  _T_5637_re = _RAND_10856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10857 = {1{`RANDOM}};
  _T_5637_im = _RAND_10857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10858 = {1{`RANDOM}};
  _T_5638_re = _RAND_10858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10859 = {1{`RANDOM}};
  _T_5638_im = _RAND_10859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10860 = {1{`RANDOM}};
  _T_5639_re = _RAND_10860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10861 = {1{`RANDOM}};
  _T_5639_im = _RAND_10861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10862 = {1{`RANDOM}};
  _T_5640_re = _RAND_10862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10863 = {1{`RANDOM}};
  _T_5640_im = _RAND_10863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10864 = {1{`RANDOM}};
  _T_5641_re = _RAND_10864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10865 = {1{`RANDOM}};
  _T_5641_im = _RAND_10865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10866 = {1{`RANDOM}};
  _T_5642_re = _RAND_10866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10867 = {1{`RANDOM}};
  _T_5642_im = _RAND_10867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10868 = {1{`RANDOM}};
  _T_5643_re = _RAND_10868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10869 = {1{`RANDOM}};
  _T_5643_im = _RAND_10869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10870 = {1{`RANDOM}};
  _T_5644_re = _RAND_10870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10871 = {1{`RANDOM}};
  _T_5644_im = _RAND_10871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10872 = {1{`RANDOM}};
  _T_5645_re = _RAND_10872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10873 = {1{`RANDOM}};
  _T_5645_im = _RAND_10873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10874 = {1{`RANDOM}};
  _T_5646_re = _RAND_10874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10875 = {1{`RANDOM}};
  _T_5646_im = _RAND_10875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10876 = {1{`RANDOM}};
  _T_5647_re = _RAND_10876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10877 = {1{`RANDOM}};
  _T_5647_im = _RAND_10877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10878 = {1{`RANDOM}};
  _T_5648_re = _RAND_10878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10879 = {1{`RANDOM}};
  _T_5648_im = _RAND_10879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10880 = {1{`RANDOM}};
  _T_5649_re = _RAND_10880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10881 = {1{`RANDOM}};
  _T_5649_im = _RAND_10881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10882 = {1{`RANDOM}};
  _T_5650_re = _RAND_10882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10883 = {1{`RANDOM}};
  _T_5650_im = _RAND_10883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10884 = {1{`RANDOM}};
  _T_5651_re = _RAND_10884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10885 = {1{`RANDOM}};
  _T_5651_im = _RAND_10885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10886 = {1{`RANDOM}};
  _T_5652_re = _RAND_10886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10887 = {1{`RANDOM}};
  _T_5652_im = _RAND_10887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10888 = {1{`RANDOM}};
  _T_5653_re = _RAND_10888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10889 = {1{`RANDOM}};
  _T_5653_im = _RAND_10889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10890 = {1{`RANDOM}};
  _T_5654_re = _RAND_10890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10891 = {1{`RANDOM}};
  _T_5654_im = _RAND_10891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10892 = {1{`RANDOM}};
  _T_5655_re = _RAND_10892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10893 = {1{`RANDOM}};
  _T_5655_im = _RAND_10893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10894 = {1{`RANDOM}};
  _T_5656_re = _RAND_10894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10895 = {1{`RANDOM}};
  _T_5656_im = _RAND_10895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10896 = {1{`RANDOM}};
  _T_5657_re = _RAND_10896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10897 = {1{`RANDOM}};
  _T_5657_im = _RAND_10897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10898 = {1{`RANDOM}};
  _T_5658_re = _RAND_10898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10899 = {1{`RANDOM}};
  _T_5658_im = _RAND_10899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10900 = {1{`RANDOM}};
  _T_5659_re = _RAND_10900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10901 = {1{`RANDOM}};
  _T_5659_im = _RAND_10901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10902 = {1{`RANDOM}};
  _T_5660_re = _RAND_10902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10903 = {1{`RANDOM}};
  _T_5660_im = _RAND_10903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10904 = {1{`RANDOM}};
  _T_5661_re = _RAND_10904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10905 = {1{`RANDOM}};
  _T_5661_im = _RAND_10905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10906 = {1{`RANDOM}};
  _T_5662_re = _RAND_10906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10907 = {1{`RANDOM}};
  _T_5662_im = _RAND_10907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10908 = {1{`RANDOM}};
  _T_5663_re = _RAND_10908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10909 = {1{`RANDOM}};
  _T_5663_im = _RAND_10909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10910 = {1{`RANDOM}};
  _T_5664_re = _RAND_10910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10911 = {1{`RANDOM}};
  _T_5664_im = _RAND_10911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10912 = {1{`RANDOM}};
  _T_5665_re = _RAND_10912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10913 = {1{`RANDOM}};
  _T_5665_im = _RAND_10913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10914 = {1{`RANDOM}};
  _T_5666_re = _RAND_10914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10915 = {1{`RANDOM}};
  _T_5666_im = _RAND_10915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10916 = {1{`RANDOM}};
  _T_5667_re = _RAND_10916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10917 = {1{`RANDOM}};
  _T_5667_im = _RAND_10917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10918 = {1{`RANDOM}};
  _T_5668_re = _RAND_10918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10919 = {1{`RANDOM}};
  _T_5668_im = _RAND_10919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10920 = {1{`RANDOM}};
  _T_5669_re = _RAND_10920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10921 = {1{`RANDOM}};
  _T_5669_im = _RAND_10921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10922 = {1{`RANDOM}};
  _T_5670_re = _RAND_10922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10923 = {1{`RANDOM}};
  _T_5670_im = _RAND_10923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10924 = {1{`RANDOM}};
  _T_5671_re = _RAND_10924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10925 = {1{`RANDOM}};
  _T_5671_im = _RAND_10925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10926 = {1{`RANDOM}};
  _T_5672_re = _RAND_10926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10927 = {1{`RANDOM}};
  _T_5672_im = _RAND_10927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10928 = {1{`RANDOM}};
  _T_5673_re = _RAND_10928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10929 = {1{`RANDOM}};
  _T_5673_im = _RAND_10929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10930 = {1{`RANDOM}};
  _T_5674_re = _RAND_10930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10931 = {1{`RANDOM}};
  _T_5674_im = _RAND_10931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10932 = {1{`RANDOM}};
  _T_5675_re = _RAND_10932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10933 = {1{`RANDOM}};
  _T_5675_im = _RAND_10933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10934 = {1{`RANDOM}};
  _T_5676_re = _RAND_10934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10935 = {1{`RANDOM}};
  _T_5676_im = _RAND_10935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10936 = {1{`RANDOM}};
  _T_5677_re = _RAND_10936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10937 = {1{`RANDOM}};
  _T_5677_im = _RAND_10937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10938 = {1{`RANDOM}};
  _T_5678_re = _RAND_10938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10939 = {1{`RANDOM}};
  _T_5678_im = _RAND_10939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10940 = {1{`RANDOM}};
  _T_5679_re = _RAND_10940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10941 = {1{`RANDOM}};
  _T_5679_im = _RAND_10941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10942 = {1{`RANDOM}};
  _T_5680_re = _RAND_10942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10943 = {1{`RANDOM}};
  _T_5680_im = _RAND_10943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10944 = {1{`RANDOM}};
  _T_5681_re = _RAND_10944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10945 = {1{`RANDOM}};
  _T_5681_im = _RAND_10945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10946 = {1{`RANDOM}};
  _T_5682_re = _RAND_10946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10947 = {1{`RANDOM}};
  _T_5682_im = _RAND_10947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10948 = {1{`RANDOM}};
  _T_5683_re = _RAND_10948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10949 = {1{`RANDOM}};
  _T_5683_im = _RAND_10949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10950 = {1{`RANDOM}};
  _T_5684_re = _RAND_10950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10951 = {1{`RANDOM}};
  _T_5684_im = _RAND_10951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10952 = {1{`RANDOM}};
  _T_5685_re = _RAND_10952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10953 = {1{`RANDOM}};
  _T_5685_im = _RAND_10953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10954 = {1{`RANDOM}};
  _T_5686_re = _RAND_10954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10955 = {1{`RANDOM}};
  _T_5686_im = _RAND_10955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10956 = {1{`RANDOM}};
  _T_5687_re = _RAND_10956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10957 = {1{`RANDOM}};
  _T_5687_im = _RAND_10957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10958 = {1{`RANDOM}};
  _T_5688_re = _RAND_10958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10959 = {1{`RANDOM}};
  _T_5688_im = _RAND_10959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10960 = {1{`RANDOM}};
  _T_5689_re = _RAND_10960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10961 = {1{`RANDOM}};
  _T_5689_im = _RAND_10961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10962 = {1{`RANDOM}};
  _T_5690_re = _RAND_10962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10963 = {1{`RANDOM}};
  _T_5690_im = _RAND_10963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10964 = {1{`RANDOM}};
  _T_5691_re = _RAND_10964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10965 = {1{`RANDOM}};
  _T_5691_im = _RAND_10965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10966 = {1{`RANDOM}};
  _T_5692_re = _RAND_10966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10967 = {1{`RANDOM}};
  _T_5692_im = _RAND_10967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10968 = {1{`RANDOM}};
  _T_5693_re = _RAND_10968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10969 = {1{`RANDOM}};
  _T_5693_im = _RAND_10969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10970 = {1{`RANDOM}};
  _T_5694_re = _RAND_10970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10971 = {1{`RANDOM}};
  _T_5694_im = _RAND_10971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10972 = {1{`RANDOM}};
  _T_5695_re = _RAND_10972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10973 = {1{`RANDOM}};
  _T_5695_im = _RAND_10973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10974 = {1{`RANDOM}};
  _T_5696_re = _RAND_10974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10975 = {1{`RANDOM}};
  _T_5696_im = _RAND_10975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10976 = {1{`RANDOM}};
  _T_5697_re = _RAND_10976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10977 = {1{`RANDOM}};
  _T_5697_im = _RAND_10977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10978 = {1{`RANDOM}};
  _T_5698_re = _RAND_10978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10979 = {1{`RANDOM}};
  _T_5698_im = _RAND_10979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10980 = {1{`RANDOM}};
  _T_5699_re = _RAND_10980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10981 = {1{`RANDOM}};
  _T_5699_im = _RAND_10981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10982 = {1{`RANDOM}};
  _T_5700_re = _RAND_10982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10983 = {1{`RANDOM}};
  _T_5700_im = _RAND_10983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10984 = {1{`RANDOM}};
  _T_5701_re = _RAND_10984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10985 = {1{`RANDOM}};
  _T_5701_im = _RAND_10985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10986 = {1{`RANDOM}};
  _T_5702_re = _RAND_10986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10987 = {1{`RANDOM}};
  _T_5702_im = _RAND_10987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10988 = {1{`RANDOM}};
  _T_5703_re = _RAND_10988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10989 = {1{`RANDOM}};
  _T_5703_im = _RAND_10989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10990 = {1{`RANDOM}};
  _T_5704_re = _RAND_10990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10991 = {1{`RANDOM}};
  _T_5704_im = _RAND_10991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10992 = {1{`RANDOM}};
  _T_5705_re = _RAND_10992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10993 = {1{`RANDOM}};
  _T_5705_im = _RAND_10993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10994 = {1{`RANDOM}};
  _T_5706_re = _RAND_10994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10995 = {1{`RANDOM}};
  _T_5706_im = _RAND_10995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10996 = {1{`RANDOM}};
  _T_5707_re = _RAND_10996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10997 = {1{`RANDOM}};
  _T_5707_im = _RAND_10997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10998 = {1{`RANDOM}};
  _T_5708_re = _RAND_10998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10999 = {1{`RANDOM}};
  _T_5708_im = _RAND_10999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11000 = {1{`RANDOM}};
  _T_5709_re = _RAND_11000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11001 = {1{`RANDOM}};
  _T_5709_im = _RAND_11001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11002 = {1{`RANDOM}};
  _T_5710_re = _RAND_11002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11003 = {1{`RANDOM}};
  _T_5710_im = _RAND_11003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11004 = {1{`RANDOM}};
  _T_5711_re = _RAND_11004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11005 = {1{`RANDOM}};
  _T_5711_im = _RAND_11005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11006 = {1{`RANDOM}};
  _T_5712_re = _RAND_11006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11007 = {1{`RANDOM}};
  _T_5712_im = _RAND_11007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11008 = {1{`RANDOM}};
  _T_5713_re = _RAND_11008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11009 = {1{`RANDOM}};
  _T_5713_im = _RAND_11009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11010 = {1{`RANDOM}};
  _T_5714_re = _RAND_11010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11011 = {1{`RANDOM}};
  _T_5714_im = _RAND_11011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11012 = {1{`RANDOM}};
  _T_5715_re = _RAND_11012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11013 = {1{`RANDOM}};
  _T_5715_im = _RAND_11013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11014 = {1{`RANDOM}};
  _T_5716_re = _RAND_11014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11015 = {1{`RANDOM}};
  _T_5716_im = _RAND_11015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11016 = {1{`RANDOM}};
  _T_5717_re = _RAND_11016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11017 = {1{`RANDOM}};
  _T_5717_im = _RAND_11017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11018 = {1{`RANDOM}};
  _T_5718_re = _RAND_11018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11019 = {1{`RANDOM}};
  _T_5718_im = _RAND_11019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11020 = {1{`RANDOM}};
  _T_5719_re = _RAND_11020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11021 = {1{`RANDOM}};
  _T_5719_im = _RAND_11021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11022 = {1{`RANDOM}};
  _T_5720_re = _RAND_11022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11023 = {1{`RANDOM}};
  _T_5720_im = _RAND_11023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11024 = {1{`RANDOM}};
  _T_5721_re = _RAND_11024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11025 = {1{`RANDOM}};
  _T_5721_im = _RAND_11025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11026 = {1{`RANDOM}};
  _T_5722_re = _RAND_11026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11027 = {1{`RANDOM}};
  _T_5722_im = _RAND_11027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11028 = {1{`RANDOM}};
  _T_5723_re = _RAND_11028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11029 = {1{`RANDOM}};
  _T_5723_im = _RAND_11029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11030 = {1{`RANDOM}};
  _T_5724_re = _RAND_11030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11031 = {1{`RANDOM}};
  _T_5724_im = _RAND_11031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11032 = {1{`RANDOM}};
  _T_5725_re = _RAND_11032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11033 = {1{`RANDOM}};
  _T_5725_im = _RAND_11033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11034 = {1{`RANDOM}};
  _T_5726_re = _RAND_11034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11035 = {1{`RANDOM}};
  _T_5726_im = _RAND_11035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11036 = {1{`RANDOM}};
  _T_5727_re = _RAND_11036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11037 = {1{`RANDOM}};
  _T_5727_im = _RAND_11037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11038 = {1{`RANDOM}};
  _T_5728_re = _RAND_11038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11039 = {1{`RANDOM}};
  _T_5728_im = _RAND_11039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11040 = {1{`RANDOM}};
  _T_5729_re = _RAND_11040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11041 = {1{`RANDOM}};
  _T_5729_im = _RAND_11041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11042 = {1{`RANDOM}};
  _T_5730_re = _RAND_11042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11043 = {1{`RANDOM}};
  _T_5730_im = _RAND_11043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11044 = {1{`RANDOM}};
  _T_5731_re = _RAND_11044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11045 = {1{`RANDOM}};
  _T_5731_im = _RAND_11045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11046 = {1{`RANDOM}};
  _T_5732_re = _RAND_11046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11047 = {1{`RANDOM}};
  _T_5732_im = _RAND_11047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11048 = {1{`RANDOM}};
  _T_5733_re = _RAND_11048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11049 = {1{`RANDOM}};
  _T_5733_im = _RAND_11049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11050 = {1{`RANDOM}};
  _T_5734_re = _RAND_11050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11051 = {1{`RANDOM}};
  _T_5734_im = _RAND_11051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11052 = {1{`RANDOM}};
  _T_5735_re = _RAND_11052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11053 = {1{`RANDOM}};
  _T_5735_im = _RAND_11053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11054 = {1{`RANDOM}};
  _T_5736_re = _RAND_11054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11055 = {1{`RANDOM}};
  _T_5736_im = _RAND_11055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11056 = {1{`RANDOM}};
  _T_5737_re = _RAND_11056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11057 = {1{`RANDOM}};
  _T_5737_im = _RAND_11057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11058 = {1{`RANDOM}};
  _T_5738_re = _RAND_11058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11059 = {1{`RANDOM}};
  _T_5738_im = _RAND_11059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11060 = {1{`RANDOM}};
  _T_5739_re = _RAND_11060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11061 = {1{`RANDOM}};
  _T_5739_im = _RAND_11061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11062 = {1{`RANDOM}};
  _T_5740_re = _RAND_11062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11063 = {1{`RANDOM}};
  _T_5740_im = _RAND_11063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11064 = {1{`RANDOM}};
  _T_5741_re = _RAND_11064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11065 = {1{`RANDOM}};
  _T_5741_im = _RAND_11065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11066 = {1{`RANDOM}};
  _T_5742_re = _RAND_11066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11067 = {1{`RANDOM}};
  _T_5742_im = _RAND_11067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11068 = {1{`RANDOM}};
  _T_5743_re = _RAND_11068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11069 = {1{`RANDOM}};
  _T_5743_im = _RAND_11069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11070 = {1{`RANDOM}};
  _T_5744_re = _RAND_11070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11071 = {1{`RANDOM}};
  _T_5744_im = _RAND_11071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11072 = {1{`RANDOM}};
  _T_5745_re = _RAND_11072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11073 = {1{`RANDOM}};
  _T_5745_im = _RAND_11073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11074 = {1{`RANDOM}};
  _T_5746_re = _RAND_11074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11075 = {1{`RANDOM}};
  _T_5746_im = _RAND_11075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11076 = {1{`RANDOM}};
  _T_5747_re = _RAND_11076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11077 = {1{`RANDOM}};
  _T_5747_im = _RAND_11077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11078 = {1{`RANDOM}};
  _T_5748_re = _RAND_11078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11079 = {1{`RANDOM}};
  _T_5748_im = _RAND_11079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11080 = {1{`RANDOM}};
  _T_5749_re = _RAND_11080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11081 = {1{`RANDOM}};
  _T_5749_im = _RAND_11081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11082 = {1{`RANDOM}};
  _T_5750_re = _RAND_11082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11083 = {1{`RANDOM}};
  _T_5750_im = _RAND_11083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11084 = {1{`RANDOM}};
  _T_5751_re = _RAND_11084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11085 = {1{`RANDOM}};
  _T_5751_im = _RAND_11085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11086 = {1{`RANDOM}};
  _T_5752_re = _RAND_11086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11087 = {1{`RANDOM}};
  _T_5752_im = _RAND_11087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11088 = {1{`RANDOM}};
  _T_5753_re = _RAND_11088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11089 = {1{`RANDOM}};
  _T_5753_im = _RAND_11089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11090 = {1{`RANDOM}};
  _T_5754_re = _RAND_11090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11091 = {1{`RANDOM}};
  _T_5754_im = _RAND_11091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11092 = {1{`RANDOM}};
  _T_5755_re = _RAND_11092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11093 = {1{`RANDOM}};
  _T_5755_im = _RAND_11093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11094 = {1{`RANDOM}};
  _T_5756_re = _RAND_11094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11095 = {1{`RANDOM}};
  _T_5756_im = _RAND_11095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11096 = {1{`RANDOM}};
  _T_5757_re = _RAND_11096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11097 = {1{`RANDOM}};
  _T_5757_im = _RAND_11097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11098 = {1{`RANDOM}};
  _T_5758_re = _RAND_11098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11099 = {1{`RANDOM}};
  _T_5758_im = _RAND_11099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11100 = {1{`RANDOM}};
  _T_5759_re = _RAND_11100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11101 = {1{`RANDOM}};
  _T_5759_im = _RAND_11101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11102 = {1{`RANDOM}};
  _T_5760_re = _RAND_11102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11103 = {1{`RANDOM}};
  _T_5760_im = _RAND_11103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11104 = {1{`RANDOM}};
  _T_5761_re = _RAND_11104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11105 = {1{`RANDOM}};
  _T_5761_im = _RAND_11105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11106 = {1{`RANDOM}};
  _T_5762_re = _RAND_11106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11107 = {1{`RANDOM}};
  _T_5762_im = _RAND_11107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11108 = {1{`RANDOM}};
  _T_5763_re = _RAND_11108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11109 = {1{`RANDOM}};
  _T_5763_im = _RAND_11109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11110 = {1{`RANDOM}};
  _T_5764_re = _RAND_11110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11111 = {1{`RANDOM}};
  _T_5764_im = _RAND_11111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11112 = {1{`RANDOM}};
  _T_5765_re = _RAND_11112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11113 = {1{`RANDOM}};
  _T_5765_im = _RAND_11113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11114 = {1{`RANDOM}};
  _T_5766_re = _RAND_11114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11115 = {1{`RANDOM}};
  _T_5766_im = _RAND_11115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11116 = {1{`RANDOM}};
  _T_5767_re = _RAND_11116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11117 = {1{`RANDOM}};
  _T_5767_im = _RAND_11117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11118 = {1{`RANDOM}};
  _T_5768_re = _RAND_11118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11119 = {1{`RANDOM}};
  _T_5768_im = _RAND_11119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11120 = {1{`RANDOM}};
  _T_5769_re = _RAND_11120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11121 = {1{`RANDOM}};
  _T_5769_im = _RAND_11121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11122 = {1{`RANDOM}};
  _T_5770_re = _RAND_11122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11123 = {1{`RANDOM}};
  _T_5770_im = _RAND_11123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11124 = {1{`RANDOM}};
  _T_5771_re = _RAND_11124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11125 = {1{`RANDOM}};
  _T_5771_im = _RAND_11125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11126 = {1{`RANDOM}};
  _T_5772_re = _RAND_11126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11127 = {1{`RANDOM}};
  _T_5772_im = _RAND_11127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11128 = {1{`RANDOM}};
  _T_5773_re = _RAND_11128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11129 = {1{`RANDOM}};
  _T_5773_im = _RAND_11129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11130 = {1{`RANDOM}};
  _T_5774_re = _RAND_11130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11131 = {1{`RANDOM}};
  _T_5774_im = _RAND_11131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11132 = {1{`RANDOM}};
  _T_5775_re = _RAND_11132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11133 = {1{`RANDOM}};
  _T_5775_im = _RAND_11133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11134 = {1{`RANDOM}};
  _T_5776_re = _RAND_11134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11135 = {1{`RANDOM}};
  _T_5776_im = _RAND_11135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11136 = {1{`RANDOM}};
  _T_5777_re = _RAND_11136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11137 = {1{`RANDOM}};
  _T_5777_im = _RAND_11137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11138 = {1{`RANDOM}};
  _T_5778_re = _RAND_11138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11139 = {1{`RANDOM}};
  _T_5778_im = _RAND_11139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11140 = {1{`RANDOM}};
  _T_5779_re = _RAND_11140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11141 = {1{`RANDOM}};
  _T_5779_im = _RAND_11141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11142 = {1{`RANDOM}};
  _T_5780_re = _RAND_11142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11143 = {1{`RANDOM}};
  _T_5780_im = _RAND_11143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11144 = {1{`RANDOM}};
  _T_5781_re = _RAND_11144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11145 = {1{`RANDOM}};
  _T_5781_im = _RAND_11145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11146 = {1{`RANDOM}};
  _T_5782_re = _RAND_11146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11147 = {1{`RANDOM}};
  _T_5782_im = _RAND_11147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11148 = {1{`RANDOM}};
  _T_5783_re = _RAND_11148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11149 = {1{`RANDOM}};
  _T_5783_im = _RAND_11149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11150 = {1{`RANDOM}};
  _T_5784_re = _RAND_11150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11151 = {1{`RANDOM}};
  _T_5784_im = _RAND_11151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11152 = {1{`RANDOM}};
  _T_5785_re = _RAND_11152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11153 = {1{`RANDOM}};
  _T_5785_im = _RAND_11153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11154 = {1{`RANDOM}};
  _T_5786_re = _RAND_11154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11155 = {1{`RANDOM}};
  _T_5786_im = _RAND_11155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11156 = {1{`RANDOM}};
  _T_5787_re = _RAND_11156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11157 = {1{`RANDOM}};
  _T_5787_im = _RAND_11157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11158 = {1{`RANDOM}};
  _T_5788_re = _RAND_11158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11159 = {1{`RANDOM}};
  _T_5788_im = _RAND_11159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11160 = {1{`RANDOM}};
  _T_5789_re = _RAND_11160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11161 = {1{`RANDOM}};
  _T_5789_im = _RAND_11161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11162 = {1{`RANDOM}};
  _T_5790_re = _RAND_11162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11163 = {1{`RANDOM}};
  _T_5790_im = _RAND_11163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11164 = {1{`RANDOM}};
  _T_5791_re = _RAND_11164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11165 = {1{`RANDOM}};
  _T_5791_im = _RAND_11165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11166 = {1{`RANDOM}};
  _T_5792_re = _RAND_11166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11167 = {1{`RANDOM}};
  _T_5792_im = _RAND_11167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11168 = {1{`RANDOM}};
  _T_5793_re = _RAND_11168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11169 = {1{`RANDOM}};
  _T_5793_im = _RAND_11169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11170 = {1{`RANDOM}};
  _T_5794_re = _RAND_11170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11171 = {1{`RANDOM}};
  _T_5794_im = _RAND_11171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11172 = {1{`RANDOM}};
  _T_5795_re = _RAND_11172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11173 = {1{`RANDOM}};
  _T_5795_im = _RAND_11173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11174 = {1{`RANDOM}};
  _T_5796_re = _RAND_11174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11175 = {1{`RANDOM}};
  _T_5796_im = _RAND_11175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11176 = {1{`RANDOM}};
  _T_5797_re = _RAND_11176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11177 = {1{`RANDOM}};
  _T_5797_im = _RAND_11177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11178 = {1{`RANDOM}};
  _T_5798_re = _RAND_11178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11179 = {1{`RANDOM}};
  _T_5798_im = _RAND_11179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11180 = {1{`RANDOM}};
  _T_5799_re = _RAND_11180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11181 = {1{`RANDOM}};
  _T_5799_im = _RAND_11181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11182 = {1{`RANDOM}};
  _T_5800_re = _RAND_11182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11183 = {1{`RANDOM}};
  _T_5800_im = _RAND_11183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11184 = {1{`RANDOM}};
  _T_5801_re = _RAND_11184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11185 = {1{`RANDOM}};
  _T_5801_im = _RAND_11185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11186 = {1{`RANDOM}};
  _T_5802_re = _RAND_11186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11187 = {1{`RANDOM}};
  _T_5802_im = _RAND_11187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11188 = {1{`RANDOM}};
  _T_5803_re = _RAND_11188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11189 = {1{`RANDOM}};
  _T_5803_im = _RAND_11189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11190 = {1{`RANDOM}};
  _T_5804_re = _RAND_11190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11191 = {1{`RANDOM}};
  _T_5804_im = _RAND_11191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11192 = {1{`RANDOM}};
  _T_5805_re = _RAND_11192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11193 = {1{`RANDOM}};
  _T_5805_im = _RAND_11193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11194 = {1{`RANDOM}};
  _T_5806_re = _RAND_11194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11195 = {1{`RANDOM}};
  _T_5806_im = _RAND_11195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11196 = {1{`RANDOM}};
  _T_5807_re = _RAND_11196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11197 = {1{`RANDOM}};
  _T_5807_im = _RAND_11197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11198 = {1{`RANDOM}};
  _T_5808_re = _RAND_11198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11199 = {1{`RANDOM}};
  _T_5808_im = _RAND_11199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11200 = {1{`RANDOM}};
  _T_5809_re = _RAND_11200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11201 = {1{`RANDOM}};
  _T_5809_im = _RAND_11201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11202 = {1{`RANDOM}};
  _T_5810_re = _RAND_11202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11203 = {1{`RANDOM}};
  _T_5810_im = _RAND_11203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11204 = {1{`RANDOM}};
  _T_5811_re = _RAND_11204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11205 = {1{`RANDOM}};
  _T_5811_im = _RAND_11205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11206 = {1{`RANDOM}};
  _T_5812_re = _RAND_11206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11207 = {1{`RANDOM}};
  _T_5812_im = _RAND_11207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11208 = {1{`RANDOM}};
  _T_5813_re = _RAND_11208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11209 = {1{`RANDOM}};
  _T_5813_im = _RAND_11209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11210 = {1{`RANDOM}};
  _T_5814_re = _RAND_11210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11211 = {1{`RANDOM}};
  _T_5814_im = _RAND_11211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11212 = {1{`RANDOM}};
  _T_5815_re = _RAND_11212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11213 = {1{`RANDOM}};
  _T_5815_im = _RAND_11213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11214 = {1{`RANDOM}};
  _T_5816_re = _RAND_11214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11215 = {1{`RANDOM}};
  _T_5816_im = _RAND_11215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11216 = {1{`RANDOM}};
  _T_5817_re = _RAND_11216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11217 = {1{`RANDOM}};
  _T_5817_im = _RAND_11217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11218 = {1{`RANDOM}};
  _T_5818_re = _RAND_11218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11219 = {1{`RANDOM}};
  _T_5818_im = _RAND_11219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11220 = {1{`RANDOM}};
  _T_5819_re = _RAND_11220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11221 = {1{`RANDOM}};
  _T_5819_im = _RAND_11221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11222 = {1{`RANDOM}};
  _T_5820_re = _RAND_11222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11223 = {1{`RANDOM}};
  _T_5820_im = _RAND_11223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11224 = {1{`RANDOM}};
  _T_5821_re = _RAND_11224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11225 = {1{`RANDOM}};
  _T_5821_im = _RAND_11225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11226 = {1{`RANDOM}};
  _T_5822_re = _RAND_11226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11227 = {1{`RANDOM}};
  _T_5822_im = _RAND_11227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11228 = {1{`RANDOM}};
  _T_5823_re = _RAND_11228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11229 = {1{`RANDOM}};
  _T_5823_im = _RAND_11229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11230 = {1{`RANDOM}};
  _T_5824_re = _RAND_11230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11231 = {1{`RANDOM}};
  _T_5824_im = _RAND_11231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11232 = {1{`RANDOM}};
  _T_5825_re = _RAND_11232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11233 = {1{`RANDOM}};
  _T_5825_im = _RAND_11233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11234 = {1{`RANDOM}};
  _T_5826_re = _RAND_11234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11235 = {1{`RANDOM}};
  _T_5826_im = _RAND_11235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11236 = {1{`RANDOM}};
  _T_5827_re = _RAND_11236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11237 = {1{`RANDOM}};
  _T_5827_im = _RAND_11237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11238 = {1{`RANDOM}};
  _T_5828_re = _RAND_11238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11239 = {1{`RANDOM}};
  _T_5828_im = _RAND_11239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11240 = {1{`RANDOM}};
  _T_5829_re = _RAND_11240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11241 = {1{`RANDOM}};
  _T_5829_im = _RAND_11241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11242 = {1{`RANDOM}};
  _T_5830_re = _RAND_11242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11243 = {1{`RANDOM}};
  _T_5830_im = _RAND_11243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11244 = {1{`RANDOM}};
  _T_5831_re = _RAND_11244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11245 = {1{`RANDOM}};
  _T_5831_im = _RAND_11245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11246 = {1{`RANDOM}};
  _T_5832_re = _RAND_11246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11247 = {1{`RANDOM}};
  _T_5832_im = _RAND_11247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11248 = {1{`RANDOM}};
  _T_5833_re = _RAND_11248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11249 = {1{`RANDOM}};
  _T_5833_im = _RAND_11249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11250 = {1{`RANDOM}};
  _T_5834_re = _RAND_11250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11251 = {1{`RANDOM}};
  _T_5834_im = _RAND_11251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11252 = {1{`RANDOM}};
  _T_5835_re = _RAND_11252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11253 = {1{`RANDOM}};
  _T_5835_im = _RAND_11253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11254 = {1{`RANDOM}};
  _T_5836_re = _RAND_11254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11255 = {1{`RANDOM}};
  _T_5836_im = _RAND_11255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11256 = {1{`RANDOM}};
  _T_5837_re = _RAND_11256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11257 = {1{`RANDOM}};
  _T_5837_im = _RAND_11257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11258 = {1{`RANDOM}};
  _T_5838_re = _RAND_11258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11259 = {1{`RANDOM}};
  _T_5838_im = _RAND_11259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11260 = {1{`RANDOM}};
  _T_5839_re = _RAND_11260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11261 = {1{`RANDOM}};
  _T_5839_im = _RAND_11261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11262 = {1{`RANDOM}};
  _T_5840_re = _RAND_11262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11263 = {1{`RANDOM}};
  _T_5840_im = _RAND_11263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11264 = {1{`RANDOM}};
  _T_5841_re = _RAND_11264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11265 = {1{`RANDOM}};
  _T_5841_im = _RAND_11265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11266 = {1{`RANDOM}};
  _T_5844_re = _RAND_11266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11267 = {1{`RANDOM}};
  _T_5844_im = _RAND_11267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11268 = {1{`RANDOM}};
  _T_5845_re = _RAND_11268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11269 = {1{`RANDOM}};
  _T_5845_im = _RAND_11269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11270 = {1{`RANDOM}};
  _T_5846_re = _RAND_11270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11271 = {1{`RANDOM}};
  _T_5846_im = _RAND_11271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11272 = {1{`RANDOM}};
  _T_5847_re = _RAND_11272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11273 = {1{`RANDOM}};
  _T_5847_im = _RAND_11273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11274 = {1{`RANDOM}};
  _T_5848_re = _RAND_11274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11275 = {1{`RANDOM}};
  _T_5848_im = _RAND_11275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11276 = {1{`RANDOM}};
  _T_5849_re = _RAND_11276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11277 = {1{`RANDOM}};
  _T_5849_im = _RAND_11277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11278 = {1{`RANDOM}};
  _T_5850_re = _RAND_11278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11279 = {1{`RANDOM}};
  _T_5850_im = _RAND_11279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11280 = {1{`RANDOM}};
  _T_5851_re = _RAND_11280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11281 = {1{`RANDOM}};
  _T_5851_im = _RAND_11281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11282 = {1{`RANDOM}};
  _T_5852_re = _RAND_11282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11283 = {1{`RANDOM}};
  _T_5852_im = _RAND_11283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11284 = {1{`RANDOM}};
  _T_5853_re = _RAND_11284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11285 = {1{`RANDOM}};
  _T_5853_im = _RAND_11285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11286 = {1{`RANDOM}};
  _T_5854_re = _RAND_11286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11287 = {1{`RANDOM}};
  _T_5854_im = _RAND_11287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11288 = {1{`RANDOM}};
  _T_5855_re = _RAND_11288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11289 = {1{`RANDOM}};
  _T_5855_im = _RAND_11289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11290 = {1{`RANDOM}};
  _T_5856_re = _RAND_11290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11291 = {1{`RANDOM}};
  _T_5856_im = _RAND_11291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11292 = {1{`RANDOM}};
  _T_5857_re = _RAND_11292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11293 = {1{`RANDOM}};
  _T_5857_im = _RAND_11293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11294 = {1{`RANDOM}};
  _T_5858_re = _RAND_11294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11295 = {1{`RANDOM}};
  _T_5858_im = _RAND_11295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11296 = {1{`RANDOM}};
  _T_5859_re = _RAND_11296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11297 = {1{`RANDOM}};
  _T_5859_im = _RAND_11297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11298 = {1{`RANDOM}};
  _T_5860_re = _RAND_11298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11299 = {1{`RANDOM}};
  _T_5860_im = _RAND_11299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11300 = {1{`RANDOM}};
  _T_5861_re = _RAND_11300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11301 = {1{`RANDOM}};
  _T_5861_im = _RAND_11301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11302 = {1{`RANDOM}};
  _T_5862_re = _RAND_11302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11303 = {1{`RANDOM}};
  _T_5862_im = _RAND_11303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11304 = {1{`RANDOM}};
  _T_5863_re = _RAND_11304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11305 = {1{`RANDOM}};
  _T_5863_im = _RAND_11305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11306 = {1{`RANDOM}};
  _T_5864_re = _RAND_11306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11307 = {1{`RANDOM}};
  _T_5864_im = _RAND_11307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11308 = {1{`RANDOM}};
  _T_5865_re = _RAND_11308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11309 = {1{`RANDOM}};
  _T_5865_im = _RAND_11309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11310 = {1{`RANDOM}};
  _T_5866_re = _RAND_11310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11311 = {1{`RANDOM}};
  _T_5866_im = _RAND_11311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11312 = {1{`RANDOM}};
  _T_5867_re = _RAND_11312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11313 = {1{`RANDOM}};
  _T_5867_im = _RAND_11313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11314 = {1{`RANDOM}};
  _T_5868_re = _RAND_11314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11315 = {1{`RANDOM}};
  _T_5868_im = _RAND_11315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11316 = {1{`RANDOM}};
  _T_5869_re = _RAND_11316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11317 = {1{`RANDOM}};
  _T_5869_im = _RAND_11317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11318 = {1{`RANDOM}};
  _T_5870_re = _RAND_11318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11319 = {1{`RANDOM}};
  _T_5870_im = _RAND_11319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11320 = {1{`RANDOM}};
  _T_5871_re = _RAND_11320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11321 = {1{`RANDOM}};
  _T_5871_im = _RAND_11321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11322 = {1{`RANDOM}};
  _T_5872_re = _RAND_11322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11323 = {1{`RANDOM}};
  _T_5872_im = _RAND_11323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11324 = {1{`RANDOM}};
  _T_5873_re = _RAND_11324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11325 = {1{`RANDOM}};
  _T_5873_im = _RAND_11325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11326 = {1{`RANDOM}};
  _T_5874_re = _RAND_11326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11327 = {1{`RANDOM}};
  _T_5874_im = _RAND_11327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11328 = {1{`RANDOM}};
  _T_5875_re = _RAND_11328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11329 = {1{`RANDOM}};
  _T_5875_im = _RAND_11329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11330 = {1{`RANDOM}};
  _T_5876_re = _RAND_11330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11331 = {1{`RANDOM}};
  _T_5876_im = _RAND_11331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11332 = {1{`RANDOM}};
  _T_5877_re = _RAND_11332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11333 = {1{`RANDOM}};
  _T_5877_im = _RAND_11333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11334 = {1{`RANDOM}};
  _T_5878_re = _RAND_11334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11335 = {1{`RANDOM}};
  _T_5878_im = _RAND_11335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11336 = {1{`RANDOM}};
  _T_5879_re = _RAND_11336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11337 = {1{`RANDOM}};
  _T_5879_im = _RAND_11337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11338 = {1{`RANDOM}};
  _T_5880_re = _RAND_11338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11339 = {1{`RANDOM}};
  _T_5880_im = _RAND_11339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11340 = {1{`RANDOM}};
  _T_5881_re = _RAND_11340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11341 = {1{`RANDOM}};
  _T_5881_im = _RAND_11341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11342 = {1{`RANDOM}};
  _T_5882_re = _RAND_11342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11343 = {1{`RANDOM}};
  _T_5882_im = _RAND_11343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11344 = {1{`RANDOM}};
  _T_5883_re = _RAND_11344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11345 = {1{`RANDOM}};
  _T_5883_im = _RAND_11345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11346 = {1{`RANDOM}};
  _T_5884_re = _RAND_11346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11347 = {1{`RANDOM}};
  _T_5884_im = _RAND_11347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11348 = {1{`RANDOM}};
  _T_5885_re = _RAND_11348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11349 = {1{`RANDOM}};
  _T_5885_im = _RAND_11349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11350 = {1{`RANDOM}};
  _T_5886_re = _RAND_11350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11351 = {1{`RANDOM}};
  _T_5886_im = _RAND_11351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11352 = {1{`RANDOM}};
  _T_5887_re = _RAND_11352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11353 = {1{`RANDOM}};
  _T_5887_im = _RAND_11353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11354 = {1{`RANDOM}};
  _T_5888_re = _RAND_11354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11355 = {1{`RANDOM}};
  _T_5888_im = _RAND_11355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11356 = {1{`RANDOM}};
  _T_5889_re = _RAND_11356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11357 = {1{`RANDOM}};
  _T_5889_im = _RAND_11357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11358 = {1{`RANDOM}};
  _T_5890_re = _RAND_11358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11359 = {1{`RANDOM}};
  _T_5890_im = _RAND_11359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11360 = {1{`RANDOM}};
  _T_5891_re = _RAND_11360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11361 = {1{`RANDOM}};
  _T_5891_im = _RAND_11361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11362 = {1{`RANDOM}};
  _T_5892_re = _RAND_11362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11363 = {1{`RANDOM}};
  _T_5892_im = _RAND_11363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11364 = {1{`RANDOM}};
  _T_5893_re = _RAND_11364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11365 = {1{`RANDOM}};
  _T_5893_im = _RAND_11365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11366 = {1{`RANDOM}};
  _T_5894_re = _RAND_11366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11367 = {1{`RANDOM}};
  _T_5894_im = _RAND_11367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11368 = {1{`RANDOM}};
  _T_5895_re = _RAND_11368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11369 = {1{`RANDOM}};
  _T_5895_im = _RAND_11369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11370 = {1{`RANDOM}};
  _T_5896_re = _RAND_11370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11371 = {1{`RANDOM}};
  _T_5896_im = _RAND_11371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11372 = {1{`RANDOM}};
  _T_5897_re = _RAND_11372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11373 = {1{`RANDOM}};
  _T_5897_im = _RAND_11373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11374 = {1{`RANDOM}};
  _T_5898_re = _RAND_11374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11375 = {1{`RANDOM}};
  _T_5898_im = _RAND_11375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11376 = {1{`RANDOM}};
  _T_5899_re = _RAND_11376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11377 = {1{`RANDOM}};
  _T_5899_im = _RAND_11377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11378 = {1{`RANDOM}};
  _T_5900_re = _RAND_11378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11379 = {1{`RANDOM}};
  _T_5900_im = _RAND_11379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11380 = {1{`RANDOM}};
  _T_5901_re = _RAND_11380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11381 = {1{`RANDOM}};
  _T_5901_im = _RAND_11381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11382 = {1{`RANDOM}};
  _T_5902_re = _RAND_11382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11383 = {1{`RANDOM}};
  _T_5902_im = _RAND_11383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11384 = {1{`RANDOM}};
  _T_5903_re = _RAND_11384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11385 = {1{`RANDOM}};
  _T_5903_im = _RAND_11385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11386 = {1{`RANDOM}};
  _T_5904_re = _RAND_11386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11387 = {1{`RANDOM}};
  _T_5904_im = _RAND_11387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11388 = {1{`RANDOM}};
  _T_5905_re = _RAND_11388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11389 = {1{`RANDOM}};
  _T_5905_im = _RAND_11389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11390 = {1{`RANDOM}};
  _T_5906_re = _RAND_11390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11391 = {1{`RANDOM}};
  _T_5906_im = _RAND_11391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11392 = {1{`RANDOM}};
  _T_5907_re = _RAND_11392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11393 = {1{`RANDOM}};
  _T_5907_im = _RAND_11393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11394 = {1{`RANDOM}};
  _T_5908_re = _RAND_11394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11395 = {1{`RANDOM}};
  _T_5908_im = _RAND_11395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11396 = {1{`RANDOM}};
  _T_5909_re = _RAND_11396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11397 = {1{`RANDOM}};
  _T_5909_im = _RAND_11397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11398 = {1{`RANDOM}};
  _T_5910_re = _RAND_11398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11399 = {1{`RANDOM}};
  _T_5910_im = _RAND_11399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11400 = {1{`RANDOM}};
  _T_5911_re = _RAND_11400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11401 = {1{`RANDOM}};
  _T_5911_im = _RAND_11401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11402 = {1{`RANDOM}};
  _T_5912_re = _RAND_11402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11403 = {1{`RANDOM}};
  _T_5912_im = _RAND_11403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11404 = {1{`RANDOM}};
  _T_5913_re = _RAND_11404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11405 = {1{`RANDOM}};
  _T_5913_im = _RAND_11405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11406 = {1{`RANDOM}};
  _T_5914_re = _RAND_11406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11407 = {1{`RANDOM}};
  _T_5914_im = _RAND_11407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11408 = {1{`RANDOM}};
  _T_5915_re = _RAND_11408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11409 = {1{`RANDOM}};
  _T_5915_im = _RAND_11409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11410 = {1{`RANDOM}};
  _T_5916_re = _RAND_11410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11411 = {1{`RANDOM}};
  _T_5916_im = _RAND_11411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11412 = {1{`RANDOM}};
  _T_5917_re = _RAND_11412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11413 = {1{`RANDOM}};
  _T_5917_im = _RAND_11413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11414 = {1{`RANDOM}};
  _T_5918_re = _RAND_11414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11415 = {1{`RANDOM}};
  _T_5918_im = _RAND_11415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11416 = {1{`RANDOM}};
  _T_5919_re = _RAND_11416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11417 = {1{`RANDOM}};
  _T_5919_im = _RAND_11417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11418 = {1{`RANDOM}};
  _T_5920_re = _RAND_11418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11419 = {1{`RANDOM}};
  _T_5920_im = _RAND_11419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11420 = {1{`RANDOM}};
  _T_5921_re = _RAND_11420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11421 = {1{`RANDOM}};
  _T_5921_im = _RAND_11421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11422 = {1{`RANDOM}};
  _T_5922_re = _RAND_11422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11423 = {1{`RANDOM}};
  _T_5922_im = _RAND_11423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11424 = {1{`RANDOM}};
  _T_5923_re = _RAND_11424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11425 = {1{`RANDOM}};
  _T_5923_im = _RAND_11425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11426 = {1{`RANDOM}};
  _T_5924_re = _RAND_11426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11427 = {1{`RANDOM}};
  _T_5924_im = _RAND_11427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11428 = {1{`RANDOM}};
  _T_5925_re = _RAND_11428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11429 = {1{`RANDOM}};
  _T_5925_im = _RAND_11429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11430 = {1{`RANDOM}};
  _T_5926_re = _RAND_11430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11431 = {1{`RANDOM}};
  _T_5926_im = _RAND_11431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11432 = {1{`RANDOM}};
  _T_5927_re = _RAND_11432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11433 = {1{`RANDOM}};
  _T_5927_im = _RAND_11433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11434 = {1{`RANDOM}};
  _T_5928_re = _RAND_11434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11435 = {1{`RANDOM}};
  _T_5928_im = _RAND_11435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11436 = {1{`RANDOM}};
  _T_5929_re = _RAND_11436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11437 = {1{`RANDOM}};
  _T_5929_im = _RAND_11437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11438 = {1{`RANDOM}};
  _T_5930_re = _RAND_11438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11439 = {1{`RANDOM}};
  _T_5930_im = _RAND_11439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11440 = {1{`RANDOM}};
  _T_5931_re = _RAND_11440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11441 = {1{`RANDOM}};
  _T_5931_im = _RAND_11441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11442 = {1{`RANDOM}};
  _T_5932_re = _RAND_11442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11443 = {1{`RANDOM}};
  _T_5932_im = _RAND_11443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11444 = {1{`RANDOM}};
  _T_5933_re = _RAND_11444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11445 = {1{`RANDOM}};
  _T_5933_im = _RAND_11445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11446 = {1{`RANDOM}};
  _T_5934_re = _RAND_11446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11447 = {1{`RANDOM}};
  _T_5934_im = _RAND_11447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11448 = {1{`RANDOM}};
  _T_5935_re = _RAND_11448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11449 = {1{`RANDOM}};
  _T_5935_im = _RAND_11449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11450 = {1{`RANDOM}};
  _T_5936_re = _RAND_11450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11451 = {1{`RANDOM}};
  _T_5936_im = _RAND_11451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11452 = {1{`RANDOM}};
  _T_5937_re = _RAND_11452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11453 = {1{`RANDOM}};
  _T_5937_im = _RAND_11453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11454 = {1{`RANDOM}};
  _T_5938_re = _RAND_11454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11455 = {1{`RANDOM}};
  _T_5938_im = _RAND_11455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11456 = {1{`RANDOM}};
  _T_5939_re = _RAND_11456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11457 = {1{`RANDOM}};
  _T_5939_im = _RAND_11457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11458 = {1{`RANDOM}};
  _T_5940_re = _RAND_11458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11459 = {1{`RANDOM}};
  _T_5940_im = _RAND_11459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11460 = {1{`RANDOM}};
  _T_5941_re = _RAND_11460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11461 = {1{`RANDOM}};
  _T_5941_im = _RAND_11461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11462 = {1{`RANDOM}};
  _T_5942_re = _RAND_11462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11463 = {1{`RANDOM}};
  _T_5942_im = _RAND_11463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11464 = {1{`RANDOM}};
  _T_5943_re = _RAND_11464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11465 = {1{`RANDOM}};
  _T_5943_im = _RAND_11465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11466 = {1{`RANDOM}};
  _T_5944_re = _RAND_11466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11467 = {1{`RANDOM}};
  _T_5944_im = _RAND_11467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11468 = {1{`RANDOM}};
  _T_5945_re = _RAND_11468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11469 = {1{`RANDOM}};
  _T_5945_im = _RAND_11469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11470 = {1{`RANDOM}};
  _T_5946_re = _RAND_11470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11471 = {1{`RANDOM}};
  _T_5946_im = _RAND_11471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11472 = {1{`RANDOM}};
  _T_5947_re = _RAND_11472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11473 = {1{`RANDOM}};
  _T_5947_im = _RAND_11473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11474 = {1{`RANDOM}};
  _T_5948_re = _RAND_11474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11475 = {1{`RANDOM}};
  _T_5948_im = _RAND_11475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11476 = {1{`RANDOM}};
  _T_5949_re = _RAND_11476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11477 = {1{`RANDOM}};
  _T_5949_im = _RAND_11477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11478 = {1{`RANDOM}};
  _T_5950_re = _RAND_11478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11479 = {1{`RANDOM}};
  _T_5950_im = _RAND_11479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11480 = {1{`RANDOM}};
  _T_5951_re = _RAND_11480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11481 = {1{`RANDOM}};
  _T_5951_im = _RAND_11481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11482 = {1{`RANDOM}};
  _T_5952_re = _RAND_11482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11483 = {1{`RANDOM}};
  _T_5952_im = _RAND_11483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11484 = {1{`RANDOM}};
  _T_5953_re = _RAND_11484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11485 = {1{`RANDOM}};
  _T_5953_im = _RAND_11485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11486 = {1{`RANDOM}};
  _T_5954_re = _RAND_11486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11487 = {1{`RANDOM}};
  _T_5954_im = _RAND_11487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11488 = {1{`RANDOM}};
  _T_5955_re = _RAND_11488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11489 = {1{`RANDOM}};
  _T_5955_im = _RAND_11489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11490 = {1{`RANDOM}};
  _T_5956_re = _RAND_11490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11491 = {1{`RANDOM}};
  _T_5956_im = _RAND_11491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11492 = {1{`RANDOM}};
  _T_5957_re = _RAND_11492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11493 = {1{`RANDOM}};
  _T_5957_im = _RAND_11493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11494 = {1{`RANDOM}};
  _T_5958_re = _RAND_11494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11495 = {1{`RANDOM}};
  _T_5958_im = _RAND_11495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11496 = {1{`RANDOM}};
  _T_5959_re = _RAND_11496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11497 = {1{`RANDOM}};
  _T_5959_im = _RAND_11497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11498 = {1{`RANDOM}};
  _T_5960_re = _RAND_11498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11499 = {1{`RANDOM}};
  _T_5960_im = _RAND_11499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11500 = {1{`RANDOM}};
  _T_5961_re = _RAND_11500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11501 = {1{`RANDOM}};
  _T_5961_im = _RAND_11501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11502 = {1{`RANDOM}};
  _T_5962_re = _RAND_11502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11503 = {1{`RANDOM}};
  _T_5962_im = _RAND_11503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11504 = {1{`RANDOM}};
  _T_5963_re = _RAND_11504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11505 = {1{`RANDOM}};
  _T_5963_im = _RAND_11505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11506 = {1{`RANDOM}};
  _T_5964_re = _RAND_11506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11507 = {1{`RANDOM}};
  _T_5964_im = _RAND_11507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11508 = {1{`RANDOM}};
  _T_5965_re = _RAND_11508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11509 = {1{`RANDOM}};
  _T_5965_im = _RAND_11509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11510 = {1{`RANDOM}};
  _T_5966_re = _RAND_11510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11511 = {1{`RANDOM}};
  _T_5966_im = _RAND_11511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11512 = {1{`RANDOM}};
  _T_5967_re = _RAND_11512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11513 = {1{`RANDOM}};
  _T_5967_im = _RAND_11513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11514 = {1{`RANDOM}};
  _T_5968_re = _RAND_11514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11515 = {1{`RANDOM}};
  _T_5968_im = _RAND_11515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11516 = {1{`RANDOM}};
  _T_5969_re = _RAND_11516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11517 = {1{`RANDOM}};
  _T_5969_im = _RAND_11517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11518 = {1{`RANDOM}};
  _T_5970_re = _RAND_11518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11519 = {1{`RANDOM}};
  _T_5970_im = _RAND_11519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11520 = {1{`RANDOM}};
  _T_5971_re = _RAND_11520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11521 = {1{`RANDOM}};
  _T_5971_im = _RAND_11521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11522 = {1{`RANDOM}};
  _T_5977_re = _RAND_11522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11523 = {1{`RANDOM}};
  _T_5977_im = _RAND_11523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11524 = {1{`RANDOM}};
  _T_5978_re = _RAND_11524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11525 = {1{`RANDOM}};
  _T_5978_im = _RAND_11525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11526 = {1{`RANDOM}};
  _T_5979_re = _RAND_11526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11527 = {1{`RANDOM}};
  _T_5979_im = _RAND_11527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11528 = {1{`RANDOM}};
  _T_5980_re = _RAND_11528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11529 = {1{`RANDOM}};
  _T_5980_im = _RAND_11529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11530 = {1{`RANDOM}};
  _T_5981_re = _RAND_11530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11531 = {1{`RANDOM}};
  _T_5981_im = _RAND_11531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11532 = {1{`RANDOM}};
  _T_5982_re = _RAND_11532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11533 = {1{`RANDOM}};
  _T_5982_im = _RAND_11533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11534 = {1{`RANDOM}};
  _T_5983_re = _RAND_11534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11535 = {1{`RANDOM}};
  _T_5983_im = _RAND_11535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11536 = {1{`RANDOM}};
  _T_5984_re = _RAND_11536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11537 = {1{`RANDOM}};
  _T_5984_im = _RAND_11537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11538 = {1{`RANDOM}};
  _T_5985_re = _RAND_11538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11539 = {1{`RANDOM}};
  _T_5985_im = _RAND_11539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11540 = {1{`RANDOM}};
  _T_5986_re = _RAND_11540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11541 = {1{`RANDOM}};
  _T_5986_im = _RAND_11541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11542 = {1{`RANDOM}};
  _T_5987_re = _RAND_11542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11543 = {1{`RANDOM}};
  _T_5987_im = _RAND_11543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11544 = {1{`RANDOM}};
  _T_5988_re = _RAND_11544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11545 = {1{`RANDOM}};
  _T_5988_im = _RAND_11545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11546 = {1{`RANDOM}};
  _T_5989_re = _RAND_11546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11547 = {1{`RANDOM}};
  _T_5989_im = _RAND_11547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11548 = {1{`RANDOM}};
  _T_5990_re = _RAND_11548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11549 = {1{`RANDOM}};
  _T_5990_im = _RAND_11549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11550 = {1{`RANDOM}};
  _T_5991_re = _RAND_11550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11551 = {1{`RANDOM}};
  _T_5991_im = _RAND_11551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11552 = {1{`RANDOM}};
  _T_5992_re = _RAND_11552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11553 = {1{`RANDOM}};
  _T_5992_im = _RAND_11553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11554 = {1{`RANDOM}};
  _T_5993_re = _RAND_11554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11555 = {1{`RANDOM}};
  _T_5993_im = _RAND_11555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11556 = {1{`RANDOM}};
  _T_5994_re = _RAND_11556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11557 = {1{`RANDOM}};
  _T_5994_im = _RAND_11557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11558 = {1{`RANDOM}};
  _T_5995_re = _RAND_11558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11559 = {1{`RANDOM}};
  _T_5995_im = _RAND_11559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11560 = {1{`RANDOM}};
  _T_5996_re = _RAND_11560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11561 = {1{`RANDOM}};
  _T_5996_im = _RAND_11561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11562 = {1{`RANDOM}};
  _T_5997_re = _RAND_11562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11563 = {1{`RANDOM}};
  _T_5997_im = _RAND_11563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11564 = {1{`RANDOM}};
  _T_5998_re = _RAND_11564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11565 = {1{`RANDOM}};
  _T_5998_im = _RAND_11565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11566 = {1{`RANDOM}};
  _T_5999_re = _RAND_11566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11567 = {1{`RANDOM}};
  _T_5999_im = _RAND_11567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11568 = {1{`RANDOM}};
  _T_6000_re = _RAND_11568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11569 = {1{`RANDOM}};
  _T_6000_im = _RAND_11569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11570 = {1{`RANDOM}};
  _T_6001_re = _RAND_11570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11571 = {1{`RANDOM}};
  _T_6001_im = _RAND_11571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11572 = {1{`RANDOM}};
  _T_6002_re = _RAND_11572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11573 = {1{`RANDOM}};
  _T_6002_im = _RAND_11573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11574 = {1{`RANDOM}};
  _T_6003_re = _RAND_11574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11575 = {1{`RANDOM}};
  _T_6003_im = _RAND_11575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11576 = {1{`RANDOM}};
  _T_6004_re = _RAND_11576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11577 = {1{`RANDOM}};
  _T_6004_im = _RAND_11577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11578 = {1{`RANDOM}};
  _T_6005_re = _RAND_11578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11579 = {1{`RANDOM}};
  _T_6005_im = _RAND_11579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11580 = {1{`RANDOM}};
  _T_6006_re = _RAND_11580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11581 = {1{`RANDOM}};
  _T_6006_im = _RAND_11581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11582 = {1{`RANDOM}};
  _T_6007_re = _RAND_11582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11583 = {1{`RANDOM}};
  _T_6007_im = _RAND_11583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11584 = {1{`RANDOM}};
  _T_6008_re = _RAND_11584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11585 = {1{`RANDOM}};
  _T_6008_im = _RAND_11585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11586 = {1{`RANDOM}};
  _T_6009_re = _RAND_11586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11587 = {1{`RANDOM}};
  _T_6009_im = _RAND_11587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11588 = {1{`RANDOM}};
  _T_6010_re = _RAND_11588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11589 = {1{`RANDOM}};
  _T_6010_im = _RAND_11589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11590 = {1{`RANDOM}};
  _T_6011_re = _RAND_11590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11591 = {1{`RANDOM}};
  _T_6011_im = _RAND_11591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11592 = {1{`RANDOM}};
  _T_6012_re = _RAND_11592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11593 = {1{`RANDOM}};
  _T_6012_im = _RAND_11593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11594 = {1{`RANDOM}};
  _T_6013_re = _RAND_11594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11595 = {1{`RANDOM}};
  _T_6013_im = _RAND_11595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11596 = {1{`RANDOM}};
  _T_6014_re = _RAND_11596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11597 = {1{`RANDOM}};
  _T_6014_im = _RAND_11597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11598 = {1{`RANDOM}};
  _T_6015_re = _RAND_11598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11599 = {1{`RANDOM}};
  _T_6015_im = _RAND_11599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11600 = {1{`RANDOM}};
  _T_6016_re = _RAND_11600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11601 = {1{`RANDOM}};
  _T_6016_im = _RAND_11601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11602 = {1{`RANDOM}};
  _T_6017_re = _RAND_11602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11603 = {1{`RANDOM}};
  _T_6017_im = _RAND_11603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11604 = {1{`RANDOM}};
  _T_6018_re = _RAND_11604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11605 = {1{`RANDOM}};
  _T_6018_im = _RAND_11605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11606 = {1{`RANDOM}};
  _T_6019_re = _RAND_11606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11607 = {1{`RANDOM}};
  _T_6019_im = _RAND_11607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11608 = {1{`RANDOM}};
  _T_6020_re = _RAND_11608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11609 = {1{`RANDOM}};
  _T_6020_im = _RAND_11609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11610 = {1{`RANDOM}};
  _T_6021_re = _RAND_11610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11611 = {1{`RANDOM}};
  _T_6021_im = _RAND_11611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11612 = {1{`RANDOM}};
  _T_6022_re = _RAND_11612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11613 = {1{`RANDOM}};
  _T_6022_im = _RAND_11613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11614 = {1{`RANDOM}};
  _T_6023_re = _RAND_11614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11615 = {1{`RANDOM}};
  _T_6023_im = _RAND_11615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11616 = {1{`RANDOM}};
  _T_6024_re = _RAND_11616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11617 = {1{`RANDOM}};
  _T_6024_im = _RAND_11617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11618 = {1{`RANDOM}};
  _T_6025_re = _RAND_11618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11619 = {1{`RANDOM}};
  _T_6025_im = _RAND_11619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11620 = {1{`RANDOM}};
  _T_6026_re = _RAND_11620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11621 = {1{`RANDOM}};
  _T_6026_im = _RAND_11621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11622 = {1{`RANDOM}};
  _T_6027_re = _RAND_11622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11623 = {1{`RANDOM}};
  _T_6027_im = _RAND_11623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11624 = {1{`RANDOM}};
  _T_6028_re = _RAND_11624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11625 = {1{`RANDOM}};
  _T_6028_im = _RAND_11625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11626 = {1{`RANDOM}};
  _T_6029_re = _RAND_11626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11627 = {1{`RANDOM}};
  _T_6029_im = _RAND_11627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11628 = {1{`RANDOM}};
  _T_6030_re = _RAND_11628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11629 = {1{`RANDOM}};
  _T_6030_im = _RAND_11629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11630 = {1{`RANDOM}};
  _T_6031_re = _RAND_11630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11631 = {1{`RANDOM}};
  _T_6031_im = _RAND_11631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11632 = {1{`RANDOM}};
  _T_6032_re = _RAND_11632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11633 = {1{`RANDOM}};
  _T_6032_im = _RAND_11633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11634 = {1{`RANDOM}};
  _T_6033_re = _RAND_11634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11635 = {1{`RANDOM}};
  _T_6033_im = _RAND_11635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11636 = {1{`RANDOM}};
  _T_6034_re = _RAND_11636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11637 = {1{`RANDOM}};
  _T_6034_im = _RAND_11637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11638 = {1{`RANDOM}};
  _T_6035_re = _RAND_11638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11639 = {1{`RANDOM}};
  _T_6035_im = _RAND_11639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11640 = {1{`RANDOM}};
  _T_6036_re = _RAND_11640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11641 = {1{`RANDOM}};
  _T_6036_im = _RAND_11641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11642 = {1{`RANDOM}};
  _T_6037_re = _RAND_11642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11643 = {1{`RANDOM}};
  _T_6037_im = _RAND_11643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11644 = {1{`RANDOM}};
  _T_6038_re = _RAND_11644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11645 = {1{`RANDOM}};
  _T_6038_im = _RAND_11645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11646 = {1{`RANDOM}};
  _T_6039_re = _RAND_11646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11647 = {1{`RANDOM}};
  _T_6039_im = _RAND_11647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11648 = {1{`RANDOM}};
  _T_6040_re = _RAND_11648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11649 = {1{`RANDOM}};
  _T_6040_im = _RAND_11649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11650 = {1{`RANDOM}};
  _T_6041_re = _RAND_11650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11651 = {1{`RANDOM}};
  _T_6041_im = _RAND_11651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11652 = {1{`RANDOM}};
  _T_6042_re = _RAND_11652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11653 = {1{`RANDOM}};
  _T_6042_im = _RAND_11653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11654 = {1{`RANDOM}};
  _T_6043_re = _RAND_11654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11655 = {1{`RANDOM}};
  _T_6043_im = _RAND_11655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11656 = {1{`RANDOM}};
  _T_6044_re = _RAND_11656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11657 = {1{`RANDOM}};
  _T_6044_im = _RAND_11657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11658 = {1{`RANDOM}};
  _T_6045_re = _RAND_11658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11659 = {1{`RANDOM}};
  _T_6045_im = _RAND_11659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11660 = {1{`RANDOM}};
  _T_6046_re = _RAND_11660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11661 = {1{`RANDOM}};
  _T_6046_im = _RAND_11661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11662 = {1{`RANDOM}};
  _T_6047_re = _RAND_11662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11663 = {1{`RANDOM}};
  _T_6047_im = _RAND_11663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11664 = {1{`RANDOM}};
  _T_6048_re = _RAND_11664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11665 = {1{`RANDOM}};
  _T_6048_im = _RAND_11665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11666 = {1{`RANDOM}};
  _T_6049_re = _RAND_11666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11667 = {1{`RANDOM}};
  _T_6049_im = _RAND_11667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11668 = {1{`RANDOM}};
  _T_6050_re = _RAND_11668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11669 = {1{`RANDOM}};
  _T_6050_im = _RAND_11669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11670 = {1{`RANDOM}};
  _T_6051_re = _RAND_11670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11671 = {1{`RANDOM}};
  _T_6051_im = _RAND_11671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11672 = {1{`RANDOM}};
  _T_6052_re = _RAND_11672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11673 = {1{`RANDOM}};
  _T_6052_im = _RAND_11673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11674 = {1{`RANDOM}};
  _T_6053_re = _RAND_11674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11675 = {1{`RANDOM}};
  _T_6053_im = _RAND_11675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11676 = {1{`RANDOM}};
  _T_6054_re = _RAND_11676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11677 = {1{`RANDOM}};
  _T_6054_im = _RAND_11677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11678 = {1{`RANDOM}};
  _T_6055_re = _RAND_11678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11679 = {1{`RANDOM}};
  _T_6055_im = _RAND_11679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11680 = {1{`RANDOM}};
  _T_6056_re = _RAND_11680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11681 = {1{`RANDOM}};
  _T_6056_im = _RAND_11681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11682 = {1{`RANDOM}};
  _T_6057_re = _RAND_11682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11683 = {1{`RANDOM}};
  _T_6057_im = _RAND_11683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11684 = {1{`RANDOM}};
  _T_6058_re = _RAND_11684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11685 = {1{`RANDOM}};
  _T_6058_im = _RAND_11685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11686 = {1{`RANDOM}};
  _T_6059_re = _RAND_11686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11687 = {1{`RANDOM}};
  _T_6059_im = _RAND_11687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11688 = {1{`RANDOM}};
  _T_6060_re = _RAND_11688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11689 = {1{`RANDOM}};
  _T_6060_im = _RAND_11689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11690 = {1{`RANDOM}};
  _T_6061_re = _RAND_11690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11691 = {1{`RANDOM}};
  _T_6061_im = _RAND_11691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11692 = {1{`RANDOM}};
  _T_6062_re = _RAND_11692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11693 = {1{`RANDOM}};
  _T_6062_im = _RAND_11693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11694 = {1{`RANDOM}};
  _T_6063_re = _RAND_11694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11695 = {1{`RANDOM}};
  _T_6063_im = _RAND_11695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11696 = {1{`RANDOM}};
  _T_6064_re = _RAND_11696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11697 = {1{`RANDOM}};
  _T_6064_im = _RAND_11697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11698 = {1{`RANDOM}};
  _T_6065_re = _RAND_11698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11699 = {1{`RANDOM}};
  _T_6065_im = _RAND_11699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11700 = {1{`RANDOM}};
  _T_6066_re = _RAND_11700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11701 = {1{`RANDOM}};
  _T_6066_im = _RAND_11701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11702 = {1{`RANDOM}};
  _T_6067_re = _RAND_11702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11703 = {1{`RANDOM}};
  _T_6067_im = _RAND_11703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11704 = {1{`RANDOM}};
  _T_6068_re = _RAND_11704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11705 = {1{`RANDOM}};
  _T_6068_im = _RAND_11705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11706 = {1{`RANDOM}};
  _T_6069_re = _RAND_11706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11707 = {1{`RANDOM}};
  _T_6069_im = _RAND_11707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11708 = {1{`RANDOM}};
  _T_6070_re = _RAND_11708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11709 = {1{`RANDOM}};
  _T_6070_im = _RAND_11709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11710 = {1{`RANDOM}};
  _T_6071_re = _RAND_11710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11711 = {1{`RANDOM}};
  _T_6071_im = _RAND_11711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11712 = {1{`RANDOM}};
  _T_6072_re = _RAND_11712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11713 = {1{`RANDOM}};
  _T_6072_im = _RAND_11713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11714 = {1{`RANDOM}};
  _T_6073_re = _RAND_11714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11715 = {1{`RANDOM}};
  _T_6073_im = _RAND_11715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11716 = {1{`RANDOM}};
  _T_6074_re = _RAND_11716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11717 = {1{`RANDOM}};
  _T_6074_im = _RAND_11717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11718 = {1{`RANDOM}};
  _T_6075_re = _RAND_11718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11719 = {1{`RANDOM}};
  _T_6075_im = _RAND_11719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11720 = {1{`RANDOM}};
  _T_6076_re = _RAND_11720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11721 = {1{`RANDOM}};
  _T_6076_im = _RAND_11721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11722 = {1{`RANDOM}};
  _T_6077_re = _RAND_11722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11723 = {1{`RANDOM}};
  _T_6077_im = _RAND_11723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11724 = {1{`RANDOM}};
  _T_6078_re = _RAND_11724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11725 = {1{`RANDOM}};
  _T_6078_im = _RAND_11725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11726 = {1{`RANDOM}};
  _T_6079_re = _RAND_11726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11727 = {1{`RANDOM}};
  _T_6079_im = _RAND_11727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11728 = {1{`RANDOM}};
  _T_6080_re = _RAND_11728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11729 = {1{`RANDOM}};
  _T_6080_im = _RAND_11729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11730 = {1{`RANDOM}};
  _T_6081_re = _RAND_11730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11731 = {1{`RANDOM}};
  _T_6081_im = _RAND_11731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11732 = {1{`RANDOM}};
  _T_6082_re = _RAND_11732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11733 = {1{`RANDOM}};
  _T_6082_im = _RAND_11733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11734 = {1{`RANDOM}};
  _T_6083_re = _RAND_11734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11735 = {1{`RANDOM}};
  _T_6083_im = _RAND_11735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11736 = {1{`RANDOM}};
  _T_6084_re = _RAND_11736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11737 = {1{`RANDOM}};
  _T_6084_im = _RAND_11737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11738 = {1{`RANDOM}};
  _T_6085_re = _RAND_11738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11739 = {1{`RANDOM}};
  _T_6085_im = _RAND_11739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11740 = {1{`RANDOM}};
  _T_6086_re = _RAND_11740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11741 = {1{`RANDOM}};
  _T_6086_im = _RAND_11741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11742 = {1{`RANDOM}};
  _T_6087_re = _RAND_11742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11743 = {1{`RANDOM}};
  _T_6087_im = _RAND_11743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11744 = {1{`RANDOM}};
  _T_6088_re = _RAND_11744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11745 = {1{`RANDOM}};
  _T_6088_im = _RAND_11745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11746 = {1{`RANDOM}};
  _T_6089_re = _RAND_11746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11747 = {1{`RANDOM}};
  _T_6089_im = _RAND_11747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11748 = {1{`RANDOM}};
  _T_6090_re = _RAND_11748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11749 = {1{`RANDOM}};
  _T_6090_im = _RAND_11749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11750 = {1{`RANDOM}};
  _T_6091_re = _RAND_11750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11751 = {1{`RANDOM}};
  _T_6091_im = _RAND_11751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11752 = {1{`RANDOM}};
  _T_6092_re = _RAND_11752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11753 = {1{`RANDOM}};
  _T_6092_im = _RAND_11753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11754 = {1{`RANDOM}};
  _T_6093_re = _RAND_11754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11755 = {1{`RANDOM}};
  _T_6093_im = _RAND_11755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11756 = {1{`RANDOM}};
  _T_6094_re = _RAND_11756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11757 = {1{`RANDOM}};
  _T_6094_im = _RAND_11757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11758 = {1{`RANDOM}};
  _T_6095_re = _RAND_11758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11759 = {1{`RANDOM}};
  _T_6095_im = _RAND_11759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11760 = {1{`RANDOM}};
  _T_6096_re = _RAND_11760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11761 = {1{`RANDOM}};
  _T_6096_im = _RAND_11761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11762 = {1{`RANDOM}};
  _T_6097_re = _RAND_11762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11763 = {1{`RANDOM}};
  _T_6097_im = _RAND_11763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11764 = {1{`RANDOM}};
  _T_6098_re = _RAND_11764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11765 = {1{`RANDOM}};
  _T_6098_im = _RAND_11765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11766 = {1{`RANDOM}};
  _T_6099_re = _RAND_11766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11767 = {1{`RANDOM}};
  _T_6099_im = _RAND_11767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11768 = {1{`RANDOM}};
  _T_6100_re = _RAND_11768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11769 = {1{`RANDOM}};
  _T_6100_im = _RAND_11769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11770 = {1{`RANDOM}};
  _T_6101_re = _RAND_11770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11771 = {1{`RANDOM}};
  _T_6101_im = _RAND_11771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11772 = {1{`RANDOM}};
  _T_6102_re = _RAND_11772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11773 = {1{`RANDOM}};
  _T_6102_im = _RAND_11773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11774 = {1{`RANDOM}};
  _T_6103_re = _RAND_11774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11775 = {1{`RANDOM}};
  _T_6103_im = _RAND_11775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11776 = {1{`RANDOM}};
  _T_6104_re = _RAND_11776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11777 = {1{`RANDOM}};
  _T_6104_im = _RAND_11777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11778 = {1{`RANDOM}};
  _T_6107_re = _RAND_11778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11779 = {1{`RANDOM}};
  _T_6107_im = _RAND_11779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11780 = {1{`RANDOM}};
  _T_6108_re = _RAND_11780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11781 = {1{`RANDOM}};
  _T_6108_im = _RAND_11781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11782 = {1{`RANDOM}};
  _T_6109_re = _RAND_11782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11783 = {1{`RANDOM}};
  _T_6109_im = _RAND_11783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11784 = {1{`RANDOM}};
  _T_6110_re = _RAND_11784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11785 = {1{`RANDOM}};
  _T_6110_im = _RAND_11785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11786 = {1{`RANDOM}};
  _T_6111_re = _RAND_11786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11787 = {1{`RANDOM}};
  _T_6111_im = _RAND_11787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11788 = {1{`RANDOM}};
  _T_6112_re = _RAND_11788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11789 = {1{`RANDOM}};
  _T_6112_im = _RAND_11789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11790 = {1{`RANDOM}};
  _T_6113_re = _RAND_11790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11791 = {1{`RANDOM}};
  _T_6113_im = _RAND_11791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11792 = {1{`RANDOM}};
  _T_6114_re = _RAND_11792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11793 = {1{`RANDOM}};
  _T_6114_im = _RAND_11793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11794 = {1{`RANDOM}};
  _T_6115_re = _RAND_11794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11795 = {1{`RANDOM}};
  _T_6115_im = _RAND_11795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11796 = {1{`RANDOM}};
  _T_6116_re = _RAND_11796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11797 = {1{`RANDOM}};
  _T_6116_im = _RAND_11797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11798 = {1{`RANDOM}};
  _T_6117_re = _RAND_11798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11799 = {1{`RANDOM}};
  _T_6117_im = _RAND_11799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11800 = {1{`RANDOM}};
  _T_6118_re = _RAND_11800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11801 = {1{`RANDOM}};
  _T_6118_im = _RAND_11801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11802 = {1{`RANDOM}};
  _T_6119_re = _RAND_11802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11803 = {1{`RANDOM}};
  _T_6119_im = _RAND_11803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11804 = {1{`RANDOM}};
  _T_6120_re = _RAND_11804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11805 = {1{`RANDOM}};
  _T_6120_im = _RAND_11805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11806 = {1{`RANDOM}};
  _T_6121_re = _RAND_11806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11807 = {1{`RANDOM}};
  _T_6121_im = _RAND_11807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11808 = {1{`RANDOM}};
  _T_6122_re = _RAND_11808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11809 = {1{`RANDOM}};
  _T_6122_im = _RAND_11809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11810 = {1{`RANDOM}};
  _T_6123_re = _RAND_11810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11811 = {1{`RANDOM}};
  _T_6123_im = _RAND_11811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11812 = {1{`RANDOM}};
  _T_6124_re = _RAND_11812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11813 = {1{`RANDOM}};
  _T_6124_im = _RAND_11813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11814 = {1{`RANDOM}};
  _T_6125_re = _RAND_11814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11815 = {1{`RANDOM}};
  _T_6125_im = _RAND_11815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11816 = {1{`RANDOM}};
  _T_6126_re = _RAND_11816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11817 = {1{`RANDOM}};
  _T_6126_im = _RAND_11817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11818 = {1{`RANDOM}};
  _T_6127_re = _RAND_11818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11819 = {1{`RANDOM}};
  _T_6127_im = _RAND_11819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11820 = {1{`RANDOM}};
  _T_6128_re = _RAND_11820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11821 = {1{`RANDOM}};
  _T_6128_im = _RAND_11821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11822 = {1{`RANDOM}};
  _T_6129_re = _RAND_11822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11823 = {1{`RANDOM}};
  _T_6129_im = _RAND_11823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11824 = {1{`RANDOM}};
  _T_6130_re = _RAND_11824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11825 = {1{`RANDOM}};
  _T_6130_im = _RAND_11825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11826 = {1{`RANDOM}};
  _T_6131_re = _RAND_11826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11827 = {1{`RANDOM}};
  _T_6131_im = _RAND_11827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11828 = {1{`RANDOM}};
  _T_6132_re = _RAND_11828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11829 = {1{`RANDOM}};
  _T_6132_im = _RAND_11829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11830 = {1{`RANDOM}};
  _T_6133_re = _RAND_11830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11831 = {1{`RANDOM}};
  _T_6133_im = _RAND_11831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11832 = {1{`RANDOM}};
  _T_6134_re = _RAND_11832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11833 = {1{`RANDOM}};
  _T_6134_im = _RAND_11833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11834 = {1{`RANDOM}};
  _T_6135_re = _RAND_11834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11835 = {1{`RANDOM}};
  _T_6135_im = _RAND_11835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11836 = {1{`RANDOM}};
  _T_6136_re = _RAND_11836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11837 = {1{`RANDOM}};
  _T_6136_im = _RAND_11837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11838 = {1{`RANDOM}};
  _T_6137_re = _RAND_11838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11839 = {1{`RANDOM}};
  _T_6137_im = _RAND_11839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11840 = {1{`RANDOM}};
  _T_6138_re = _RAND_11840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11841 = {1{`RANDOM}};
  _T_6138_im = _RAND_11841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11842 = {1{`RANDOM}};
  _T_6139_re = _RAND_11842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11843 = {1{`RANDOM}};
  _T_6139_im = _RAND_11843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11844 = {1{`RANDOM}};
  _T_6140_re = _RAND_11844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11845 = {1{`RANDOM}};
  _T_6140_im = _RAND_11845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11846 = {1{`RANDOM}};
  _T_6141_re = _RAND_11846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11847 = {1{`RANDOM}};
  _T_6141_im = _RAND_11847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11848 = {1{`RANDOM}};
  _T_6142_re = _RAND_11848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11849 = {1{`RANDOM}};
  _T_6142_im = _RAND_11849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11850 = {1{`RANDOM}};
  _T_6143_re = _RAND_11850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11851 = {1{`RANDOM}};
  _T_6143_im = _RAND_11851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11852 = {1{`RANDOM}};
  _T_6144_re = _RAND_11852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11853 = {1{`RANDOM}};
  _T_6144_im = _RAND_11853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11854 = {1{`RANDOM}};
  _T_6145_re = _RAND_11854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11855 = {1{`RANDOM}};
  _T_6145_im = _RAND_11855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11856 = {1{`RANDOM}};
  _T_6146_re = _RAND_11856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11857 = {1{`RANDOM}};
  _T_6146_im = _RAND_11857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11858 = {1{`RANDOM}};
  _T_6147_re = _RAND_11858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11859 = {1{`RANDOM}};
  _T_6147_im = _RAND_11859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11860 = {1{`RANDOM}};
  _T_6148_re = _RAND_11860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11861 = {1{`RANDOM}};
  _T_6148_im = _RAND_11861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11862 = {1{`RANDOM}};
  _T_6149_re = _RAND_11862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11863 = {1{`RANDOM}};
  _T_6149_im = _RAND_11863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11864 = {1{`RANDOM}};
  _T_6150_re = _RAND_11864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11865 = {1{`RANDOM}};
  _T_6150_im = _RAND_11865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11866 = {1{`RANDOM}};
  _T_6151_re = _RAND_11866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11867 = {1{`RANDOM}};
  _T_6151_im = _RAND_11867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11868 = {1{`RANDOM}};
  _T_6152_re = _RAND_11868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11869 = {1{`RANDOM}};
  _T_6152_im = _RAND_11869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11870 = {1{`RANDOM}};
  _T_6153_re = _RAND_11870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11871 = {1{`RANDOM}};
  _T_6153_im = _RAND_11871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11872 = {1{`RANDOM}};
  _T_6154_re = _RAND_11872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11873 = {1{`RANDOM}};
  _T_6154_im = _RAND_11873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11874 = {1{`RANDOM}};
  _T_6155_re = _RAND_11874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11875 = {1{`RANDOM}};
  _T_6155_im = _RAND_11875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11876 = {1{`RANDOM}};
  _T_6156_re = _RAND_11876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11877 = {1{`RANDOM}};
  _T_6156_im = _RAND_11877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11878 = {1{`RANDOM}};
  _T_6157_re = _RAND_11878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11879 = {1{`RANDOM}};
  _T_6157_im = _RAND_11879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11880 = {1{`RANDOM}};
  _T_6158_re = _RAND_11880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11881 = {1{`RANDOM}};
  _T_6158_im = _RAND_11881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11882 = {1{`RANDOM}};
  _T_6159_re = _RAND_11882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11883 = {1{`RANDOM}};
  _T_6159_im = _RAND_11883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11884 = {1{`RANDOM}};
  _T_6160_re = _RAND_11884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11885 = {1{`RANDOM}};
  _T_6160_im = _RAND_11885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11886 = {1{`RANDOM}};
  _T_6161_re = _RAND_11886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11887 = {1{`RANDOM}};
  _T_6161_im = _RAND_11887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11888 = {1{`RANDOM}};
  _T_6162_re = _RAND_11888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11889 = {1{`RANDOM}};
  _T_6162_im = _RAND_11889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11890 = {1{`RANDOM}};
  _T_6163_re = _RAND_11890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11891 = {1{`RANDOM}};
  _T_6163_im = _RAND_11891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11892 = {1{`RANDOM}};
  _T_6164_re = _RAND_11892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11893 = {1{`RANDOM}};
  _T_6164_im = _RAND_11893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11894 = {1{`RANDOM}};
  _T_6165_re = _RAND_11894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11895 = {1{`RANDOM}};
  _T_6165_im = _RAND_11895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11896 = {1{`RANDOM}};
  _T_6166_re = _RAND_11896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11897 = {1{`RANDOM}};
  _T_6166_im = _RAND_11897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11898 = {1{`RANDOM}};
  _T_6167_re = _RAND_11898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11899 = {1{`RANDOM}};
  _T_6167_im = _RAND_11899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11900 = {1{`RANDOM}};
  _T_6168_re = _RAND_11900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11901 = {1{`RANDOM}};
  _T_6168_im = _RAND_11901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11902 = {1{`RANDOM}};
  _T_6169_re = _RAND_11902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11903 = {1{`RANDOM}};
  _T_6169_im = _RAND_11903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11904 = {1{`RANDOM}};
  _T_6170_re = _RAND_11904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11905 = {1{`RANDOM}};
  _T_6170_im = _RAND_11905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11906 = {1{`RANDOM}};
  _T_6176_re = _RAND_11906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11907 = {1{`RANDOM}};
  _T_6176_im = _RAND_11907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11908 = {1{`RANDOM}};
  _T_6177_re = _RAND_11908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11909 = {1{`RANDOM}};
  _T_6177_im = _RAND_11909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11910 = {1{`RANDOM}};
  _T_6178_re = _RAND_11910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11911 = {1{`RANDOM}};
  _T_6178_im = _RAND_11911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11912 = {1{`RANDOM}};
  _T_6179_re = _RAND_11912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11913 = {1{`RANDOM}};
  _T_6179_im = _RAND_11913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11914 = {1{`RANDOM}};
  _T_6180_re = _RAND_11914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11915 = {1{`RANDOM}};
  _T_6180_im = _RAND_11915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11916 = {1{`RANDOM}};
  _T_6181_re = _RAND_11916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11917 = {1{`RANDOM}};
  _T_6181_im = _RAND_11917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11918 = {1{`RANDOM}};
  _T_6182_re = _RAND_11918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11919 = {1{`RANDOM}};
  _T_6182_im = _RAND_11919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11920 = {1{`RANDOM}};
  _T_6183_re = _RAND_11920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11921 = {1{`RANDOM}};
  _T_6183_im = _RAND_11921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11922 = {1{`RANDOM}};
  _T_6184_re = _RAND_11922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11923 = {1{`RANDOM}};
  _T_6184_im = _RAND_11923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11924 = {1{`RANDOM}};
  _T_6185_re = _RAND_11924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11925 = {1{`RANDOM}};
  _T_6185_im = _RAND_11925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11926 = {1{`RANDOM}};
  _T_6186_re = _RAND_11926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11927 = {1{`RANDOM}};
  _T_6186_im = _RAND_11927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11928 = {1{`RANDOM}};
  _T_6187_re = _RAND_11928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11929 = {1{`RANDOM}};
  _T_6187_im = _RAND_11929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11930 = {1{`RANDOM}};
  _T_6188_re = _RAND_11930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11931 = {1{`RANDOM}};
  _T_6188_im = _RAND_11931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11932 = {1{`RANDOM}};
  _T_6189_re = _RAND_11932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11933 = {1{`RANDOM}};
  _T_6189_im = _RAND_11933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11934 = {1{`RANDOM}};
  _T_6190_re = _RAND_11934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11935 = {1{`RANDOM}};
  _T_6190_im = _RAND_11935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11936 = {1{`RANDOM}};
  _T_6191_re = _RAND_11936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11937 = {1{`RANDOM}};
  _T_6191_im = _RAND_11937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11938 = {1{`RANDOM}};
  _T_6192_re = _RAND_11938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11939 = {1{`RANDOM}};
  _T_6192_im = _RAND_11939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11940 = {1{`RANDOM}};
  _T_6193_re = _RAND_11940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11941 = {1{`RANDOM}};
  _T_6193_im = _RAND_11941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11942 = {1{`RANDOM}};
  _T_6194_re = _RAND_11942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11943 = {1{`RANDOM}};
  _T_6194_im = _RAND_11943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11944 = {1{`RANDOM}};
  _T_6195_re = _RAND_11944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11945 = {1{`RANDOM}};
  _T_6195_im = _RAND_11945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11946 = {1{`RANDOM}};
  _T_6196_re = _RAND_11946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11947 = {1{`RANDOM}};
  _T_6196_im = _RAND_11947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11948 = {1{`RANDOM}};
  _T_6197_re = _RAND_11948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11949 = {1{`RANDOM}};
  _T_6197_im = _RAND_11949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11950 = {1{`RANDOM}};
  _T_6198_re = _RAND_11950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11951 = {1{`RANDOM}};
  _T_6198_im = _RAND_11951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11952 = {1{`RANDOM}};
  _T_6199_re = _RAND_11952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11953 = {1{`RANDOM}};
  _T_6199_im = _RAND_11953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11954 = {1{`RANDOM}};
  _T_6200_re = _RAND_11954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11955 = {1{`RANDOM}};
  _T_6200_im = _RAND_11955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11956 = {1{`RANDOM}};
  _T_6201_re = _RAND_11956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11957 = {1{`RANDOM}};
  _T_6201_im = _RAND_11957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11958 = {1{`RANDOM}};
  _T_6202_re = _RAND_11958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11959 = {1{`RANDOM}};
  _T_6202_im = _RAND_11959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11960 = {1{`RANDOM}};
  _T_6203_re = _RAND_11960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11961 = {1{`RANDOM}};
  _T_6203_im = _RAND_11961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11962 = {1{`RANDOM}};
  _T_6204_re = _RAND_11962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11963 = {1{`RANDOM}};
  _T_6204_im = _RAND_11963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11964 = {1{`RANDOM}};
  _T_6205_re = _RAND_11964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11965 = {1{`RANDOM}};
  _T_6205_im = _RAND_11965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11966 = {1{`RANDOM}};
  _T_6206_re = _RAND_11966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11967 = {1{`RANDOM}};
  _T_6206_im = _RAND_11967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11968 = {1{`RANDOM}};
  _T_6207_re = _RAND_11968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11969 = {1{`RANDOM}};
  _T_6207_im = _RAND_11969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11970 = {1{`RANDOM}};
  _T_6208_re = _RAND_11970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11971 = {1{`RANDOM}};
  _T_6208_im = _RAND_11971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11972 = {1{`RANDOM}};
  _T_6209_re = _RAND_11972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11973 = {1{`RANDOM}};
  _T_6209_im = _RAND_11973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11974 = {1{`RANDOM}};
  _T_6210_re = _RAND_11974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11975 = {1{`RANDOM}};
  _T_6210_im = _RAND_11975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11976 = {1{`RANDOM}};
  _T_6211_re = _RAND_11976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11977 = {1{`RANDOM}};
  _T_6211_im = _RAND_11977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11978 = {1{`RANDOM}};
  _T_6212_re = _RAND_11978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11979 = {1{`RANDOM}};
  _T_6212_im = _RAND_11979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11980 = {1{`RANDOM}};
  _T_6213_re = _RAND_11980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11981 = {1{`RANDOM}};
  _T_6213_im = _RAND_11981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11982 = {1{`RANDOM}};
  _T_6214_re = _RAND_11982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11983 = {1{`RANDOM}};
  _T_6214_im = _RAND_11983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11984 = {1{`RANDOM}};
  _T_6215_re = _RAND_11984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11985 = {1{`RANDOM}};
  _T_6215_im = _RAND_11985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11986 = {1{`RANDOM}};
  _T_6216_re = _RAND_11986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11987 = {1{`RANDOM}};
  _T_6216_im = _RAND_11987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11988 = {1{`RANDOM}};
  _T_6217_re = _RAND_11988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11989 = {1{`RANDOM}};
  _T_6217_im = _RAND_11989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11990 = {1{`RANDOM}};
  _T_6218_re = _RAND_11990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11991 = {1{`RANDOM}};
  _T_6218_im = _RAND_11991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11992 = {1{`RANDOM}};
  _T_6219_re = _RAND_11992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11993 = {1{`RANDOM}};
  _T_6219_im = _RAND_11993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11994 = {1{`RANDOM}};
  _T_6220_re = _RAND_11994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11995 = {1{`RANDOM}};
  _T_6220_im = _RAND_11995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11996 = {1{`RANDOM}};
  _T_6221_re = _RAND_11996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11997 = {1{`RANDOM}};
  _T_6221_im = _RAND_11997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11998 = {1{`RANDOM}};
  _T_6222_re = _RAND_11998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11999 = {1{`RANDOM}};
  _T_6222_im = _RAND_11999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12000 = {1{`RANDOM}};
  _T_6223_re = _RAND_12000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12001 = {1{`RANDOM}};
  _T_6223_im = _RAND_12001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12002 = {1{`RANDOM}};
  _T_6224_re = _RAND_12002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12003 = {1{`RANDOM}};
  _T_6224_im = _RAND_12003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12004 = {1{`RANDOM}};
  _T_6225_re = _RAND_12004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12005 = {1{`RANDOM}};
  _T_6225_im = _RAND_12005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12006 = {1{`RANDOM}};
  _T_6226_re = _RAND_12006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12007 = {1{`RANDOM}};
  _T_6226_im = _RAND_12007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12008 = {1{`RANDOM}};
  _T_6227_re = _RAND_12008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12009 = {1{`RANDOM}};
  _T_6227_im = _RAND_12009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12010 = {1{`RANDOM}};
  _T_6228_re = _RAND_12010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12011 = {1{`RANDOM}};
  _T_6228_im = _RAND_12011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12012 = {1{`RANDOM}};
  _T_6229_re = _RAND_12012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12013 = {1{`RANDOM}};
  _T_6229_im = _RAND_12013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12014 = {1{`RANDOM}};
  _T_6230_re = _RAND_12014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12015 = {1{`RANDOM}};
  _T_6230_im = _RAND_12015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12016 = {1{`RANDOM}};
  _T_6231_re = _RAND_12016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12017 = {1{`RANDOM}};
  _T_6231_im = _RAND_12017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12018 = {1{`RANDOM}};
  _T_6232_re = _RAND_12018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12019 = {1{`RANDOM}};
  _T_6232_im = _RAND_12019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12020 = {1{`RANDOM}};
  _T_6233_re = _RAND_12020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12021 = {1{`RANDOM}};
  _T_6233_im = _RAND_12021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12022 = {1{`RANDOM}};
  _T_6234_re = _RAND_12022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12023 = {1{`RANDOM}};
  _T_6234_im = _RAND_12023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12024 = {1{`RANDOM}};
  _T_6235_re = _RAND_12024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12025 = {1{`RANDOM}};
  _T_6235_im = _RAND_12025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12026 = {1{`RANDOM}};
  _T_6236_re = _RAND_12026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12027 = {1{`RANDOM}};
  _T_6236_im = _RAND_12027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12028 = {1{`RANDOM}};
  _T_6237_re = _RAND_12028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12029 = {1{`RANDOM}};
  _T_6237_im = _RAND_12029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12030 = {1{`RANDOM}};
  _T_6238_re = _RAND_12030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12031 = {1{`RANDOM}};
  _T_6238_im = _RAND_12031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12032 = {1{`RANDOM}};
  _T_6239_re = _RAND_12032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12033 = {1{`RANDOM}};
  _T_6239_im = _RAND_12033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12034 = {1{`RANDOM}};
  _T_6242_re = _RAND_12034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12035 = {1{`RANDOM}};
  _T_6242_im = _RAND_12035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12036 = {1{`RANDOM}};
  _T_6243_re = _RAND_12036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12037 = {1{`RANDOM}};
  _T_6243_im = _RAND_12037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12038 = {1{`RANDOM}};
  _T_6244_re = _RAND_12038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12039 = {1{`RANDOM}};
  _T_6244_im = _RAND_12039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12040 = {1{`RANDOM}};
  _T_6245_re = _RAND_12040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12041 = {1{`RANDOM}};
  _T_6245_im = _RAND_12041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12042 = {1{`RANDOM}};
  _T_6246_re = _RAND_12042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12043 = {1{`RANDOM}};
  _T_6246_im = _RAND_12043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12044 = {1{`RANDOM}};
  _T_6247_re = _RAND_12044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12045 = {1{`RANDOM}};
  _T_6247_im = _RAND_12045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12046 = {1{`RANDOM}};
  _T_6248_re = _RAND_12046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12047 = {1{`RANDOM}};
  _T_6248_im = _RAND_12047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12048 = {1{`RANDOM}};
  _T_6249_re = _RAND_12048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12049 = {1{`RANDOM}};
  _T_6249_im = _RAND_12049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12050 = {1{`RANDOM}};
  _T_6250_re = _RAND_12050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12051 = {1{`RANDOM}};
  _T_6250_im = _RAND_12051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12052 = {1{`RANDOM}};
  _T_6251_re = _RAND_12052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12053 = {1{`RANDOM}};
  _T_6251_im = _RAND_12053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12054 = {1{`RANDOM}};
  _T_6252_re = _RAND_12054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12055 = {1{`RANDOM}};
  _T_6252_im = _RAND_12055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12056 = {1{`RANDOM}};
  _T_6253_re = _RAND_12056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12057 = {1{`RANDOM}};
  _T_6253_im = _RAND_12057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12058 = {1{`RANDOM}};
  _T_6254_re = _RAND_12058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12059 = {1{`RANDOM}};
  _T_6254_im = _RAND_12059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12060 = {1{`RANDOM}};
  _T_6255_re = _RAND_12060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12061 = {1{`RANDOM}};
  _T_6255_im = _RAND_12061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12062 = {1{`RANDOM}};
  _T_6256_re = _RAND_12062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12063 = {1{`RANDOM}};
  _T_6256_im = _RAND_12063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12064 = {1{`RANDOM}};
  _T_6257_re = _RAND_12064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12065 = {1{`RANDOM}};
  _T_6257_im = _RAND_12065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12066 = {1{`RANDOM}};
  _T_6258_re = _RAND_12066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12067 = {1{`RANDOM}};
  _T_6258_im = _RAND_12067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12068 = {1{`RANDOM}};
  _T_6259_re = _RAND_12068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12069 = {1{`RANDOM}};
  _T_6259_im = _RAND_12069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12070 = {1{`RANDOM}};
  _T_6260_re = _RAND_12070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12071 = {1{`RANDOM}};
  _T_6260_im = _RAND_12071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12072 = {1{`RANDOM}};
  _T_6261_re = _RAND_12072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12073 = {1{`RANDOM}};
  _T_6261_im = _RAND_12073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12074 = {1{`RANDOM}};
  _T_6262_re = _RAND_12074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12075 = {1{`RANDOM}};
  _T_6262_im = _RAND_12075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12076 = {1{`RANDOM}};
  _T_6263_re = _RAND_12076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12077 = {1{`RANDOM}};
  _T_6263_im = _RAND_12077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12078 = {1{`RANDOM}};
  _T_6264_re = _RAND_12078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12079 = {1{`RANDOM}};
  _T_6264_im = _RAND_12079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12080 = {1{`RANDOM}};
  _T_6265_re = _RAND_12080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12081 = {1{`RANDOM}};
  _T_6265_im = _RAND_12081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12082 = {1{`RANDOM}};
  _T_6266_re = _RAND_12082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12083 = {1{`RANDOM}};
  _T_6266_im = _RAND_12083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12084 = {1{`RANDOM}};
  _T_6267_re = _RAND_12084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12085 = {1{`RANDOM}};
  _T_6267_im = _RAND_12085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12086 = {1{`RANDOM}};
  _T_6268_re = _RAND_12086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12087 = {1{`RANDOM}};
  _T_6268_im = _RAND_12087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12088 = {1{`RANDOM}};
  _T_6269_re = _RAND_12088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12089 = {1{`RANDOM}};
  _T_6269_im = _RAND_12089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12090 = {1{`RANDOM}};
  _T_6270_re = _RAND_12090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12091 = {1{`RANDOM}};
  _T_6270_im = _RAND_12091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12092 = {1{`RANDOM}};
  _T_6271_re = _RAND_12092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12093 = {1{`RANDOM}};
  _T_6271_im = _RAND_12093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12094 = {1{`RANDOM}};
  _T_6272_re = _RAND_12094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12095 = {1{`RANDOM}};
  _T_6272_im = _RAND_12095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12096 = {1{`RANDOM}};
  _T_6273_re = _RAND_12096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12097 = {1{`RANDOM}};
  _T_6273_im = _RAND_12097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12098 = {1{`RANDOM}};
  _T_6279_re = _RAND_12098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12099 = {1{`RANDOM}};
  _T_6279_im = _RAND_12099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12100 = {1{`RANDOM}};
  _T_6280_re = _RAND_12100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12101 = {1{`RANDOM}};
  _T_6280_im = _RAND_12101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12102 = {1{`RANDOM}};
  _T_6281_re = _RAND_12102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12103 = {1{`RANDOM}};
  _T_6281_im = _RAND_12103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12104 = {1{`RANDOM}};
  _T_6282_re = _RAND_12104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12105 = {1{`RANDOM}};
  _T_6282_im = _RAND_12105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12106 = {1{`RANDOM}};
  _T_6283_re = _RAND_12106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12107 = {1{`RANDOM}};
  _T_6283_im = _RAND_12107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12108 = {1{`RANDOM}};
  _T_6284_re = _RAND_12108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12109 = {1{`RANDOM}};
  _T_6284_im = _RAND_12109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12110 = {1{`RANDOM}};
  _T_6285_re = _RAND_12110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12111 = {1{`RANDOM}};
  _T_6285_im = _RAND_12111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12112 = {1{`RANDOM}};
  _T_6286_re = _RAND_12112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12113 = {1{`RANDOM}};
  _T_6286_im = _RAND_12113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12114 = {1{`RANDOM}};
  _T_6287_re = _RAND_12114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12115 = {1{`RANDOM}};
  _T_6287_im = _RAND_12115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12116 = {1{`RANDOM}};
  _T_6288_re = _RAND_12116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12117 = {1{`RANDOM}};
  _T_6288_im = _RAND_12117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12118 = {1{`RANDOM}};
  _T_6289_re = _RAND_12118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12119 = {1{`RANDOM}};
  _T_6289_im = _RAND_12119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12120 = {1{`RANDOM}};
  _T_6290_re = _RAND_12120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12121 = {1{`RANDOM}};
  _T_6290_im = _RAND_12121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12122 = {1{`RANDOM}};
  _T_6291_re = _RAND_12122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12123 = {1{`RANDOM}};
  _T_6291_im = _RAND_12123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12124 = {1{`RANDOM}};
  _T_6292_re = _RAND_12124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12125 = {1{`RANDOM}};
  _T_6292_im = _RAND_12125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12126 = {1{`RANDOM}};
  _T_6293_re = _RAND_12126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12127 = {1{`RANDOM}};
  _T_6293_im = _RAND_12127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12128 = {1{`RANDOM}};
  _T_6294_re = _RAND_12128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12129 = {1{`RANDOM}};
  _T_6294_im = _RAND_12129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12130 = {1{`RANDOM}};
  _T_6295_re = _RAND_12130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12131 = {1{`RANDOM}};
  _T_6295_im = _RAND_12131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12132 = {1{`RANDOM}};
  _T_6296_re = _RAND_12132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12133 = {1{`RANDOM}};
  _T_6296_im = _RAND_12133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12134 = {1{`RANDOM}};
  _T_6297_re = _RAND_12134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12135 = {1{`RANDOM}};
  _T_6297_im = _RAND_12135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12136 = {1{`RANDOM}};
  _T_6298_re = _RAND_12136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12137 = {1{`RANDOM}};
  _T_6298_im = _RAND_12137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12138 = {1{`RANDOM}};
  _T_6299_re = _RAND_12138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12139 = {1{`RANDOM}};
  _T_6299_im = _RAND_12139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12140 = {1{`RANDOM}};
  _T_6300_re = _RAND_12140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12141 = {1{`RANDOM}};
  _T_6300_im = _RAND_12141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12142 = {1{`RANDOM}};
  _T_6301_re = _RAND_12142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12143 = {1{`RANDOM}};
  _T_6301_im = _RAND_12143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12144 = {1{`RANDOM}};
  _T_6302_re = _RAND_12144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12145 = {1{`RANDOM}};
  _T_6302_im = _RAND_12145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12146 = {1{`RANDOM}};
  _T_6303_re = _RAND_12146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12147 = {1{`RANDOM}};
  _T_6303_im = _RAND_12147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12148 = {1{`RANDOM}};
  _T_6304_re = _RAND_12148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12149 = {1{`RANDOM}};
  _T_6304_im = _RAND_12149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12150 = {1{`RANDOM}};
  _T_6305_re = _RAND_12150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12151 = {1{`RANDOM}};
  _T_6305_im = _RAND_12151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12152 = {1{`RANDOM}};
  _T_6306_re = _RAND_12152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12153 = {1{`RANDOM}};
  _T_6306_im = _RAND_12153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12154 = {1{`RANDOM}};
  _T_6307_re = _RAND_12154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12155 = {1{`RANDOM}};
  _T_6307_im = _RAND_12155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12156 = {1{`RANDOM}};
  _T_6308_re = _RAND_12156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12157 = {1{`RANDOM}};
  _T_6308_im = _RAND_12157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12158 = {1{`RANDOM}};
  _T_6309_re = _RAND_12158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12159 = {1{`RANDOM}};
  _T_6309_im = _RAND_12159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12160 = {1{`RANDOM}};
  _T_6310_re = _RAND_12160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12161 = {1{`RANDOM}};
  _T_6310_im = _RAND_12161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12162 = {1{`RANDOM}};
  _T_6313_re = _RAND_12162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12163 = {1{`RANDOM}};
  _T_6313_im = _RAND_12163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12164 = {1{`RANDOM}};
  _T_6314_re = _RAND_12164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12165 = {1{`RANDOM}};
  _T_6314_im = _RAND_12165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12166 = {1{`RANDOM}};
  _T_6315_re = _RAND_12166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12167 = {1{`RANDOM}};
  _T_6315_im = _RAND_12167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12168 = {1{`RANDOM}};
  _T_6316_re = _RAND_12168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12169 = {1{`RANDOM}};
  _T_6316_im = _RAND_12169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12170 = {1{`RANDOM}};
  _T_6317_re = _RAND_12170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12171 = {1{`RANDOM}};
  _T_6317_im = _RAND_12171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12172 = {1{`RANDOM}};
  _T_6318_re = _RAND_12172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12173 = {1{`RANDOM}};
  _T_6318_im = _RAND_12173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12174 = {1{`RANDOM}};
  _T_6319_re = _RAND_12174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12175 = {1{`RANDOM}};
  _T_6319_im = _RAND_12175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12176 = {1{`RANDOM}};
  _T_6320_re = _RAND_12176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12177 = {1{`RANDOM}};
  _T_6320_im = _RAND_12177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12178 = {1{`RANDOM}};
  _T_6321_re = _RAND_12178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12179 = {1{`RANDOM}};
  _T_6321_im = _RAND_12179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12180 = {1{`RANDOM}};
  _T_6322_re = _RAND_12180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12181 = {1{`RANDOM}};
  _T_6322_im = _RAND_12181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12182 = {1{`RANDOM}};
  _T_6323_re = _RAND_12182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12183 = {1{`RANDOM}};
  _T_6323_im = _RAND_12183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12184 = {1{`RANDOM}};
  _T_6324_re = _RAND_12184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12185 = {1{`RANDOM}};
  _T_6324_im = _RAND_12185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12186 = {1{`RANDOM}};
  _T_6325_re = _RAND_12186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12187 = {1{`RANDOM}};
  _T_6325_im = _RAND_12187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12188 = {1{`RANDOM}};
  _T_6326_re = _RAND_12188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12189 = {1{`RANDOM}};
  _T_6326_im = _RAND_12189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12190 = {1{`RANDOM}};
  _T_6327_re = _RAND_12190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12191 = {1{`RANDOM}};
  _T_6327_im = _RAND_12191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12192 = {1{`RANDOM}};
  _T_6328_re = _RAND_12192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12193 = {1{`RANDOM}};
  _T_6328_im = _RAND_12193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12194 = {1{`RANDOM}};
  _T_6334_re = _RAND_12194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12195 = {1{`RANDOM}};
  _T_6334_im = _RAND_12195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12196 = {1{`RANDOM}};
  _T_6335_re = _RAND_12196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12197 = {1{`RANDOM}};
  _T_6335_im = _RAND_12197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12198 = {1{`RANDOM}};
  _T_6336_re = _RAND_12198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12199 = {1{`RANDOM}};
  _T_6336_im = _RAND_12199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12200 = {1{`RANDOM}};
  _T_6337_re = _RAND_12200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12201 = {1{`RANDOM}};
  _T_6337_im = _RAND_12201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12202 = {1{`RANDOM}};
  _T_6338_re = _RAND_12202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12203 = {1{`RANDOM}};
  _T_6338_im = _RAND_12203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12204 = {1{`RANDOM}};
  _T_6339_re = _RAND_12204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12205 = {1{`RANDOM}};
  _T_6339_im = _RAND_12205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12206 = {1{`RANDOM}};
  _T_6340_re = _RAND_12206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12207 = {1{`RANDOM}};
  _T_6340_im = _RAND_12207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12208 = {1{`RANDOM}};
  _T_6341_re = _RAND_12208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12209 = {1{`RANDOM}};
  _T_6341_im = _RAND_12209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12210 = {1{`RANDOM}};
  _T_6342_re = _RAND_12210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12211 = {1{`RANDOM}};
  _T_6342_im = _RAND_12211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12212 = {1{`RANDOM}};
  _T_6343_re = _RAND_12212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12213 = {1{`RANDOM}};
  _T_6343_im = _RAND_12213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12214 = {1{`RANDOM}};
  _T_6344_re = _RAND_12214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12215 = {1{`RANDOM}};
  _T_6344_im = _RAND_12215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12216 = {1{`RANDOM}};
  _T_6345_re = _RAND_12216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12217 = {1{`RANDOM}};
  _T_6345_im = _RAND_12217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12218 = {1{`RANDOM}};
  _T_6346_re = _RAND_12218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12219 = {1{`RANDOM}};
  _T_6346_im = _RAND_12219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12220 = {1{`RANDOM}};
  _T_6347_re = _RAND_12220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12221 = {1{`RANDOM}};
  _T_6347_im = _RAND_12221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12222 = {1{`RANDOM}};
  _T_6348_re = _RAND_12222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12223 = {1{`RANDOM}};
  _T_6348_im = _RAND_12223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12224 = {1{`RANDOM}};
  _T_6349_re = _RAND_12224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12225 = {1{`RANDOM}};
  _T_6349_im = _RAND_12225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12226 = {1{`RANDOM}};
  _T_6352_re = _RAND_12226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12227 = {1{`RANDOM}};
  _T_6352_im = _RAND_12227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12228 = {1{`RANDOM}};
  _T_6353_re = _RAND_12228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12229 = {1{`RANDOM}};
  _T_6353_im = _RAND_12229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12230 = {1{`RANDOM}};
  _T_6354_re = _RAND_12230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12231 = {1{`RANDOM}};
  _T_6354_im = _RAND_12231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12232 = {1{`RANDOM}};
  _T_6355_re = _RAND_12232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12233 = {1{`RANDOM}};
  _T_6355_im = _RAND_12233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12234 = {1{`RANDOM}};
  _T_6356_re = _RAND_12234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12235 = {1{`RANDOM}};
  _T_6356_im = _RAND_12235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12236 = {1{`RANDOM}};
  _T_6357_re = _RAND_12236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12237 = {1{`RANDOM}};
  _T_6357_im = _RAND_12237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12238 = {1{`RANDOM}};
  _T_6358_re = _RAND_12238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12239 = {1{`RANDOM}};
  _T_6358_im = _RAND_12239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12240 = {1{`RANDOM}};
  _T_6359_re = _RAND_12240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12241 = {1{`RANDOM}};
  _T_6359_im = _RAND_12241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12242 = {1{`RANDOM}};
  _T_6365_re = _RAND_12242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12243 = {1{`RANDOM}};
  _T_6365_im = _RAND_12243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12244 = {1{`RANDOM}};
  _T_6366_re = _RAND_12244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12245 = {1{`RANDOM}};
  _T_6366_im = _RAND_12245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12246 = {1{`RANDOM}};
  _T_6367_re = _RAND_12246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12247 = {1{`RANDOM}};
  _T_6367_im = _RAND_12247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12248 = {1{`RANDOM}};
  _T_6368_re = _RAND_12248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12249 = {1{`RANDOM}};
  _T_6368_im = _RAND_12249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12250 = {1{`RANDOM}};
  _T_6369_re = _RAND_12250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12251 = {1{`RANDOM}};
  _T_6369_im = _RAND_12251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12252 = {1{`RANDOM}};
  _T_6370_re = _RAND_12252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12253 = {1{`RANDOM}};
  _T_6370_im = _RAND_12253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12254 = {1{`RANDOM}};
  _T_6371_re = _RAND_12254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12255 = {1{`RANDOM}};
  _T_6371_im = _RAND_12255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12256 = {1{`RANDOM}};
  _T_6372_re = _RAND_12256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12257 = {1{`RANDOM}};
  _T_6372_im = _RAND_12257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12258 = {1{`RANDOM}};
  _T_6375_re = _RAND_12258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12259 = {1{`RANDOM}};
  _T_6375_im = _RAND_12259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12260 = {1{`RANDOM}};
  _T_6376_re = _RAND_12260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12261 = {1{`RANDOM}};
  _T_6376_im = _RAND_12261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12262 = {1{`RANDOM}};
  _T_6377_re = _RAND_12262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12263 = {1{`RANDOM}};
  _T_6377_im = _RAND_12263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12264 = {1{`RANDOM}};
  _T_6378_re = _RAND_12264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12265 = {1{`RANDOM}};
  _T_6378_im = _RAND_12265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12266 = {1{`RANDOM}};
  _T_6384_re = _RAND_12266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12267 = {1{`RANDOM}};
  _T_6384_im = _RAND_12267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12268 = {1{`RANDOM}};
  _T_6385_re = _RAND_12268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12269 = {1{`RANDOM}};
  _T_6385_im = _RAND_12269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12270 = {1{`RANDOM}};
  _T_6386_re = _RAND_12270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12271 = {1{`RANDOM}};
  _T_6386_im = _RAND_12271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12272 = {1{`RANDOM}};
  _T_6387_re = _RAND_12272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12273 = {1{`RANDOM}};
  _T_6387_im = _RAND_12273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12274 = {1{`RANDOM}};
  _T_6390_re = _RAND_12274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12275 = {1{`RANDOM}};
  _T_6390_im = _RAND_12275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12276 = {1{`RANDOM}};
  _T_6391_re = _RAND_12276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12277 = {1{`RANDOM}};
  _T_6391_im = _RAND_12277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12278 = {1{`RANDOM}};
  _T_6397_re = _RAND_12278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12279 = {1{`RANDOM}};
  _T_6397_im = _RAND_12279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12280 = {1{`RANDOM}};
  _T_6398_re = _RAND_12280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12281 = {1{`RANDOM}};
  _T_6398_im = _RAND_12281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12282 = {1{`RANDOM}};
  _T_6401_re = _RAND_12282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12283 = {1{`RANDOM}};
  _T_6401_im = _RAND_12283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12284 = {1{`RANDOM}};
  out1D1_re = _RAND_12284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12285 = {1{`RANDOM}};
  out1D1_im = _RAND_12285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12286 = {1{`RANDOM}};
  _T_6402_re = _RAND_12286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12287 = {1{`RANDOM}};
  _T_6402_im = _RAND_12287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12288 = {1{`RANDOM}};
  _T_6403_re = _RAND_12288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12289 = {1{`RANDOM}};
  _T_6403_im = _RAND_12289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 12'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    cntD1 <= cnt;
    _T_189_re <= io_dIn_re;
    _T_189_im <= io_dIn_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_538_re <= _T_537_re;
    _T_538_im <= _T_537_im;
    _T_539_re <= _T_538_re;
    _T_539_im <= _T_538_im;
    _T_540_re <= _T_539_re;
    _T_540_im <= _T_539_im;
    _T_541_re <= _T_540_re;
    _T_541_im <= _T_540_im;
    _T_542_re <= _T_541_re;
    _T_542_im <= _T_541_im;
    _T_543_re <= _T_542_re;
    _T_543_im <= _T_542_im;
    _T_544_re <= _T_543_re;
    _T_544_im <= _T_543_im;
    _T_545_re <= _T_544_re;
    _T_545_im <= _T_544_im;
    _T_546_re <= _T_545_re;
    _T_546_im <= _T_545_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_674_re <= _T_673_re;
    _T_674_im <= _T_673_im;
    _T_675_re <= _T_674_re;
    _T_675_im <= _T_674_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_739_re <= _T_738_re;
    _T_739_im <= _T_738_im;
    _T_740_re <= _T_739_re;
    _T_740_im <= _T_739_im;
    _T_741_re <= _T_740_re;
    _T_741_im <= _T_740_im;
    _T_742_re <= _T_741_re;
    _T_742_im <= _T_741_im;
    _T_743_re <= _T_742_re;
    _T_743_im <= _T_742_im;
    _T_744_re <= _T_743_re;
    _T_744_im <= _T_743_im;
    _T_745_re <= _T_744_re;
    _T_745_im <= _T_744_im;
    _T_746_re <= _T_745_re;
    _T_746_im <= _T_745_im;
    _T_747_re <= _T_746_re;
    _T_747_im <= _T_746_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_844_re <= _T_843_re;
    _T_844_im <= _T_843_im;
    _T_845_re <= _T_844_re;
    _T_845_im <= _T_844_im;
    _T_846_re <= _T_845_re;
    _T_846_im <= _T_845_im;
    _T_847_re <= _T_846_re;
    _T_847_im <= _T_846_im;
    _T_848_re <= _T_847_re;
    _T_848_im <= _T_847_im;
    _T_849_re <= _T_848_re;
    _T_849_im <= _T_848_im;
    _T_850_re <= _T_849_re;
    _T_850_im <= _T_849_im;
    _T_851_re <= _T_850_re;
    _T_851_im <= _T_850_im;
    _T_852_re <= _T_851_re;
    _T_852_im <= _T_851_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_882_re <= _T_881_re;
    _T_882_im <= _T_881_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_884_re <= _T_883_re;
    _T_884_im <= _T_883_im;
    _T_885_re <= _T_884_re;
    _T_885_im <= _T_884_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_901_re <= _T_900_re;
    _T_901_im <= _T_900_im;
    _T_902_re <= _T_901_re;
    _T_902_im <= _T_901_im;
    _T_903_re <= _T_902_re;
    _T_903_im <= _T_902_im;
    _T_904_re <= _T_903_re;
    _T_904_im <= _T_903_im;
    _T_905_re <= _T_904_re;
    _T_905_im <= _T_904_im;
    _T_906_re <= _T_905_re;
    _T_906_im <= _T_905_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_908_re <= _T_907_re;
    _T_908_im <= _T_907_im;
    _T_909_re <= _T_908_re;
    _T_909_im <= _T_908_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_911_re <= _T_910_re;
    _T_911_im <= _T_910_im;
    _T_912_re <= _T_911_re;
    _T_912_im <= _T_911_im;
    _T_913_re <= _T_912_re;
    _T_913_im <= _T_912_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_923_re <= _T_922_re;
    _T_923_im <= _T_922_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_929_re <= _T_928_re;
    _T_929_im <= _T_928_im;
    _T_930_re <= _T_929_re;
    _T_930_im <= _T_929_im;
    _T_931_re <= _T_930_re;
    _T_931_im <= _T_930_im;
    _T_932_re <= _T_931_re;
    _T_932_im <= _T_931_im;
    _T_933_re <= _T_932_re;
    _T_933_im <= _T_932_im;
    _T_934_re <= _T_933_re;
    _T_934_im <= _T_933_im;
    _T_935_re <= _T_934_re;
    _T_935_im <= _T_934_im;
    _T_936_re <= _T_935_re;
    _T_936_im <= _T_935_im;
    _T_937_re <= _T_936_re;
    _T_937_im <= _T_936_im;
    _T_938_re <= _T_937_re;
    _T_938_im <= _T_937_im;
    _T_939_re <= _T_938_re;
    _T_939_im <= _T_938_im;
    _T_940_re <= _T_939_re;
    _T_940_im <= _T_939_im;
    _T_941_re <= _T_940_re;
    _T_941_im <= _T_940_im;
    _T_942_re <= _T_941_re;
    _T_942_im <= _T_941_im;
    _T_943_re <= _T_942_re;
    _T_943_im <= _T_942_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_947_re <= _T_946_re;
    _T_947_im <= _T_946_im;
    _T_948_re <= _T_947_re;
    _T_948_im <= _T_947_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_950_re <= _T_949_re;
    _T_950_im <= _T_949_im;
    _T_951_re <= _T_950_re;
    _T_951_im <= _T_950_im;
    _T_952_re <= _T_951_re;
    _T_952_im <= _T_951_im;
    _T_953_re <= _T_952_re;
    _T_953_im <= _T_952_im;
    _T_954_re <= _T_953_re;
    _T_954_im <= _T_953_im;
    _T_955_re <= _T_954_re;
    _T_955_im <= _T_954_im;
    _T_956_re <= _T_955_re;
    _T_956_im <= _T_955_im;
    _T_957_re <= _T_956_re;
    _T_957_im <= _T_956_im;
    _T_958_re <= _T_957_re;
    _T_958_im <= _T_957_im;
    _T_959_re <= _T_958_re;
    _T_959_im <= _T_958_im;
    _T_960_re <= _T_959_re;
    _T_960_im <= _T_959_im;
    _T_961_re <= _T_960_re;
    _T_961_im <= _T_960_im;
    _T_962_re <= _T_961_re;
    _T_962_im <= _T_961_im;
    _T_963_re <= _T_962_re;
    _T_963_im <= _T_962_im;
    _T_964_re <= _T_963_re;
    _T_964_im <= _T_963_im;
    _T_965_re <= _T_964_re;
    _T_965_im <= _T_964_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_967_re <= _T_966_re;
    _T_967_im <= _T_966_im;
    _T_968_re <= _T_967_re;
    _T_968_im <= _T_967_im;
    _T_969_re <= _T_968_re;
    _T_969_im <= _T_968_im;
    _T_970_re <= _T_969_re;
    _T_970_im <= _T_969_im;
    _T_971_re <= _T_970_re;
    _T_971_im <= _T_970_im;
    _T_972_re <= _T_971_re;
    _T_972_im <= _T_971_im;
    _T_973_re <= _T_972_re;
    _T_973_im <= _T_972_im;
    _T_974_re <= _T_973_re;
    _T_974_im <= _T_973_im;
    _T_975_re <= _T_974_re;
    _T_975_im <= _T_974_im;
    _T_976_re <= _T_975_re;
    _T_976_im <= _T_975_im;
    _T_977_re <= _T_976_re;
    _T_977_im <= _T_976_im;
    _T_978_re <= _T_977_re;
    _T_978_im <= _T_977_im;
    _T_979_re <= _T_978_re;
    _T_979_im <= _T_978_im;
    _T_980_re <= _T_979_re;
    _T_980_im <= _T_979_im;
    _T_981_re <= _T_980_re;
    _T_981_im <= _T_980_im;
    _T_982_re <= _T_981_re;
    _T_982_im <= _T_981_im;
    _T_983_re <= _T_982_re;
    _T_983_im <= _T_982_im;
    _T_984_re <= _T_983_re;
    _T_984_im <= _T_983_im;
    _T_985_re <= _T_984_re;
    _T_985_im <= _T_984_im;
    _T_986_re <= _T_985_re;
    _T_986_im <= _T_985_im;
    _T_987_re <= _T_986_re;
    _T_987_im <= _T_986_im;
    _T_988_re <= _T_987_re;
    _T_988_im <= _T_987_im;
    _T_989_re <= _T_988_re;
    _T_989_im <= _T_988_im;
    _T_990_re <= _T_989_re;
    _T_990_im <= _T_989_im;
    _T_991_re <= _T_990_re;
    _T_991_im <= _T_990_im;
    _T_992_re <= _T_991_re;
    _T_992_im <= _T_991_im;
    _T_993_re <= _T_992_re;
    _T_993_im <= _T_992_im;
    _T_994_re <= _T_993_re;
    _T_994_im <= _T_993_im;
    _T_995_re <= _T_994_re;
    _T_995_im <= _T_994_im;
    _T_996_re <= _T_995_re;
    _T_996_im <= _T_995_im;
    _T_997_re <= _T_996_re;
    _T_997_im <= _T_996_im;
    _T_998_re <= _T_997_re;
    _T_998_im <= _T_997_im;
    _T_999_re <= _T_998_re;
    _T_999_im <= _T_998_im;
    _T_1000_re <= _T_999_re;
    _T_1000_im <= _T_999_im;
    _T_1001_re <= _T_1000_re;
    _T_1001_im <= _T_1000_im;
    _T_1002_re <= _T_1001_re;
    _T_1002_im <= _T_1001_im;
    _T_1003_re <= _T_1002_re;
    _T_1003_im <= _T_1002_im;
    _T_1004_re <= _T_1003_re;
    _T_1004_im <= _T_1003_im;
    _T_1005_re <= _T_1004_re;
    _T_1005_im <= _T_1004_im;
    _T_1006_re <= _T_1005_re;
    _T_1006_im <= _T_1005_im;
    _T_1007_re <= _T_1006_re;
    _T_1007_im <= _T_1006_im;
    _T_1008_re <= _T_1007_re;
    _T_1008_im <= _T_1007_im;
    _T_1009_re <= _T_1008_re;
    _T_1009_im <= _T_1008_im;
    _T_1010_re <= _T_1009_re;
    _T_1010_im <= _T_1009_im;
    _T_1011_re <= _T_1010_re;
    _T_1011_im <= _T_1010_im;
    _T_1012_re <= _T_1011_re;
    _T_1012_im <= _T_1011_im;
    _T_1013_re <= _T_1012_re;
    _T_1013_im <= _T_1012_im;
    _T_1014_re <= _T_1013_re;
    _T_1014_im <= _T_1013_im;
    _T_1015_re <= _T_1014_re;
    _T_1015_im <= _T_1014_im;
    _T_1016_re <= _T_1015_re;
    _T_1016_im <= _T_1015_im;
    _T_1017_re <= _T_1016_re;
    _T_1017_im <= _T_1016_im;
    _T_1018_re <= _T_1017_re;
    _T_1018_im <= _T_1017_im;
    _T_1019_re <= _T_1018_re;
    _T_1019_im <= _T_1018_im;
    _T_1020_re <= _T_1019_re;
    _T_1020_im <= _T_1019_im;
    _T_1021_re <= _T_1020_re;
    _T_1021_im <= _T_1020_im;
    _T_1022_re <= _T_1021_re;
    _T_1022_im <= _T_1021_im;
    _T_1023_re <= _T_1022_re;
    _T_1023_im <= _T_1022_im;
    _T_1024_re <= _T_1023_re;
    _T_1024_im <= _T_1023_im;
    _T_1025_re <= _T_1024_re;
    _T_1025_im <= _T_1024_im;
    _T_1026_re <= _T_1025_re;
    _T_1026_im <= _T_1025_im;
    _T_1027_re <= _T_1026_re;
    _T_1027_im <= _T_1026_im;
    _T_1028_re <= _T_1027_re;
    _T_1028_im <= _T_1027_im;
    _T_1029_re <= _T_1028_re;
    _T_1029_im <= _T_1028_im;
    _T_1030_re <= _T_1029_re;
    _T_1030_im <= _T_1029_im;
    _T_1031_re <= _T_1030_re;
    _T_1031_im <= _T_1030_im;
    _T_1032_re <= _T_1031_re;
    _T_1032_im <= _T_1031_im;
    _T_1033_re <= _T_1032_re;
    _T_1033_im <= _T_1032_im;
    _T_1034_re <= _T_1033_re;
    _T_1034_im <= _T_1033_im;
    _T_1035_re <= _T_1034_re;
    _T_1035_im <= _T_1034_im;
    _T_1036_re <= _T_1035_re;
    _T_1036_im <= _T_1035_im;
    _T_1037_re <= _T_1036_re;
    _T_1037_im <= _T_1036_im;
    _T_1038_re <= _T_1037_re;
    _T_1038_im <= _T_1037_im;
    _T_1039_re <= _T_1038_re;
    _T_1039_im <= _T_1038_im;
    _T_1040_re <= _T_1039_re;
    _T_1040_im <= _T_1039_im;
    _T_1041_re <= _T_1040_re;
    _T_1041_im <= _T_1040_im;
    _T_1042_re <= _T_1041_re;
    _T_1042_im <= _T_1041_im;
    _T_1043_re <= _T_1042_re;
    _T_1043_im <= _T_1042_im;
    _T_1044_re <= _T_1043_re;
    _T_1044_im <= _T_1043_im;
    _T_1045_re <= _T_1044_re;
    _T_1045_im <= _T_1044_im;
    _T_1046_re <= _T_1045_re;
    _T_1046_im <= _T_1045_im;
    _T_1047_re <= _T_1046_re;
    _T_1047_im <= _T_1046_im;
    _T_1048_re <= _T_1047_re;
    _T_1048_im <= _T_1047_im;
    _T_1049_re <= _T_1048_re;
    _T_1049_im <= _T_1048_im;
    _T_1050_re <= _T_1049_re;
    _T_1050_im <= _T_1049_im;
    _T_1051_re <= _T_1050_re;
    _T_1051_im <= _T_1050_im;
    _T_1052_re <= _T_1051_re;
    _T_1052_im <= _T_1051_im;
    _T_1053_re <= _T_1052_re;
    _T_1053_im <= _T_1052_im;
    _T_1054_re <= _T_1053_re;
    _T_1054_im <= _T_1053_im;
    _T_1055_re <= _T_1054_re;
    _T_1055_im <= _T_1054_im;
    _T_1056_re <= _T_1055_re;
    _T_1056_im <= _T_1055_im;
    _T_1057_re <= _T_1056_re;
    _T_1057_im <= _T_1056_im;
    _T_1058_re <= _T_1057_re;
    _T_1058_im <= _T_1057_im;
    _T_1059_re <= _T_1058_re;
    _T_1059_im <= _T_1058_im;
    _T_1060_re <= _T_1059_re;
    _T_1060_im <= _T_1059_im;
    _T_1061_re <= _T_1060_re;
    _T_1061_im <= _T_1060_im;
    _T_1062_re <= _T_1061_re;
    _T_1062_im <= _T_1061_im;
    _T_1063_re <= _T_1062_re;
    _T_1063_im <= _T_1062_im;
    _T_1064_re <= _T_1063_re;
    _T_1064_im <= _T_1063_im;
    _T_1065_re <= _T_1064_re;
    _T_1065_im <= _T_1064_im;
    _T_1066_re <= _T_1065_re;
    _T_1066_im <= _T_1065_im;
    _T_1067_re <= _T_1066_re;
    _T_1067_im <= _T_1066_im;
    _T_1068_re <= _T_1067_re;
    _T_1068_im <= _T_1067_im;
    _T_1069_re <= _T_1068_re;
    _T_1069_im <= _T_1068_im;
    _T_1070_re <= _T_1069_re;
    _T_1070_im <= _T_1069_im;
    _T_1071_re <= _T_1070_re;
    _T_1071_im <= _T_1070_im;
    _T_1072_re <= _T_1071_re;
    _T_1072_im <= _T_1071_im;
    _T_1073_re <= _T_1072_re;
    _T_1073_im <= _T_1072_im;
    _T_1074_re <= _T_1073_re;
    _T_1074_im <= _T_1073_im;
    _T_1075_re <= _T_1074_re;
    _T_1075_im <= _T_1074_im;
    _T_1076_re <= _T_1075_re;
    _T_1076_im <= _T_1075_im;
    _T_1077_re <= _T_1076_re;
    _T_1077_im <= _T_1076_im;
    _T_1078_re <= _T_1077_re;
    _T_1078_im <= _T_1077_im;
    _T_1079_re <= _T_1078_re;
    _T_1079_im <= _T_1078_im;
    _T_1080_re <= _T_1079_re;
    _T_1080_im <= _T_1079_im;
    _T_1081_re <= _T_1080_re;
    _T_1081_im <= _T_1080_im;
    _T_1082_re <= _T_1081_re;
    _T_1082_im <= _T_1081_im;
    _T_1083_re <= _T_1082_re;
    _T_1083_im <= _T_1082_im;
    _T_1084_re <= _T_1083_re;
    _T_1084_im <= _T_1083_im;
    _T_1085_re <= _T_1084_re;
    _T_1085_im <= _T_1084_im;
    _T_1086_re <= _T_1085_re;
    _T_1086_im <= _T_1085_im;
    _T_1087_re <= _T_1086_re;
    _T_1087_im <= _T_1086_im;
    _T_1088_re <= _T_1087_re;
    _T_1088_im <= _T_1087_im;
    _T_1089_re <= _T_1088_re;
    _T_1089_im <= _T_1088_im;
    _T_1090_re <= _T_1089_re;
    _T_1090_im <= _T_1089_im;
    _T_1091_re <= _T_1090_re;
    _T_1091_im <= _T_1090_im;
    _T_1092_re <= _T_1091_re;
    _T_1092_im <= _T_1091_im;
    _T_1093_re <= _T_1092_re;
    _T_1093_im <= _T_1092_im;
    _T_1094_re <= _T_1093_re;
    _T_1094_im <= _T_1093_im;
    _T_1095_re <= _T_1094_re;
    _T_1095_im <= _T_1094_im;
    _T_1096_re <= _T_1095_re;
    _T_1096_im <= _T_1095_im;
    _T_1097_re <= _T_1096_re;
    _T_1097_im <= _T_1096_im;
    _T_1098_re <= _T_1097_re;
    _T_1098_im <= _T_1097_im;
    _T_1099_re <= _T_1098_re;
    _T_1099_im <= _T_1098_im;
    _T_1100_re <= _T_1099_re;
    _T_1100_im <= _T_1099_im;
    _T_1101_re <= _T_1100_re;
    _T_1101_im <= _T_1100_im;
    _T_1102_re <= _T_1101_re;
    _T_1102_im <= _T_1101_im;
    _T_1103_re <= _T_1102_re;
    _T_1103_im <= _T_1102_im;
    _T_1104_re <= _T_1103_re;
    _T_1104_im <= _T_1103_im;
    _T_1105_re <= _T_1104_re;
    _T_1105_im <= _T_1104_im;
    _T_1106_re <= _T_1105_re;
    _T_1106_im <= _T_1105_im;
    _T_1107_re <= _T_1106_re;
    _T_1107_im <= _T_1106_im;
    _T_1108_re <= _T_1107_re;
    _T_1108_im <= _T_1107_im;
    _T_1109_re <= _T_1108_re;
    _T_1109_im <= _T_1108_im;
    _T_1110_re <= _T_1109_re;
    _T_1110_im <= _T_1109_im;
    _T_1111_re <= _T_1110_re;
    _T_1111_im <= _T_1110_im;
    _T_1112_re <= _T_1111_re;
    _T_1112_im <= _T_1111_im;
    _T_1113_re <= _T_1112_re;
    _T_1113_im <= _T_1112_im;
    _T_1114_re <= _T_1113_re;
    _T_1114_im <= _T_1113_im;
    _T_1115_re <= _T_1114_re;
    _T_1115_im <= _T_1114_im;
    _T_1116_re <= _T_1115_re;
    _T_1116_im <= _T_1115_im;
    _T_1117_re <= _T_1116_re;
    _T_1117_im <= _T_1116_im;
    _T_1118_re <= _T_1117_re;
    _T_1118_im <= _T_1117_im;
    _T_1119_re <= _T_1118_re;
    _T_1119_im <= _T_1118_im;
    _T_1120_re <= _T_1119_re;
    _T_1120_im <= _T_1119_im;
    _T_1121_re <= _T_1120_re;
    _T_1121_im <= _T_1120_im;
    _T_1122_re <= _T_1121_re;
    _T_1122_im <= _T_1121_im;
    _T_1123_re <= _T_1122_re;
    _T_1123_im <= _T_1122_im;
    _T_1124_re <= _T_1123_re;
    _T_1124_im <= _T_1123_im;
    _T_1125_re <= _T_1124_re;
    _T_1125_im <= _T_1124_im;
    _T_1126_re <= _T_1125_re;
    _T_1126_im <= _T_1125_im;
    _T_1127_re <= _T_1126_re;
    _T_1127_im <= _T_1126_im;
    _T_1128_re <= _T_1127_re;
    _T_1128_im <= _T_1127_im;
    _T_1129_re <= _T_1128_re;
    _T_1129_im <= _T_1128_im;
    _T_1130_re <= _T_1129_re;
    _T_1130_im <= _T_1129_im;
    _T_1131_re <= _T_1130_re;
    _T_1131_im <= _T_1130_im;
    _T_1132_re <= _T_1131_re;
    _T_1132_im <= _T_1131_im;
    _T_1133_re <= _T_1132_re;
    _T_1133_im <= _T_1132_im;
    _T_1134_re <= _T_1133_re;
    _T_1134_im <= _T_1133_im;
    _T_1135_re <= _T_1134_re;
    _T_1135_im <= _T_1134_im;
    _T_1136_re <= _T_1135_re;
    _T_1136_im <= _T_1135_im;
    _T_1137_re <= _T_1136_re;
    _T_1137_im <= _T_1136_im;
    _T_1138_re <= _T_1137_re;
    _T_1138_im <= _T_1137_im;
    _T_1139_re <= _T_1138_re;
    _T_1139_im <= _T_1138_im;
    _T_1140_re <= _T_1139_re;
    _T_1140_im <= _T_1139_im;
    _T_1141_re <= _T_1140_re;
    _T_1141_im <= _T_1140_im;
    _T_1142_re <= _T_1141_re;
    _T_1142_im <= _T_1141_im;
    _T_1143_re <= _T_1142_re;
    _T_1143_im <= _T_1142_im;
    _T_1144_re <= _T_1143_re;
    _T_1144_im <= _T_1143_im;
    _T_1145_re <= _T_1144_re;
    _T_1145_im <= _T_1144_im;
    _T_1146_re <= _T_1145_re;
    _T_1146_im <= _T_1145_im;
    _T_1147_re <= _T_1146_re;
    _T_1147_im <= _T_1146_im;
    _T_1148_re <= _T_1147_re;
    _T_1148_im <= _T_1147_im;
    _T_1149_re <= _T_1148_re;
    _T_1149_im <= _T_1148_im;
    _T_1150_re <= _T_1149_re;
    _T_1150_im <= _T_1149_im;
    _T_1151_re <= _T_1150_re;
    _T_1151_im <= _T_1150_im;
    _T_1152_re <= _T_1151_re;
    _T_1152_im <= _T_1151_im;
    _T_1153_re <= _T_1152_re;
    _T_1153_im <= _T_1152_im;
    _T_1154_re <= _T_1153_re;
    _T_1154_im <= _T_1153_im;
    _T_1155_re <= _T_1154_re;
    _T_1155_im <= _T_1154_im;
    _T_1156_re <= _T_1155_re;
    _T_1156_im <= _T_1155_im;
    _T_1157_re <= _T_1156_re;
    _T_1157_im <= _T_1156_im;
    _T_1158_re <= _T_1157_re;
    _T_1158_im <= _T_1157_im;
    _T_1159_re <= _T_1158_re;
    _T_1159_im <= _T_1158_im;
    _T_1160_re <= _T_1159_re;
    _T_1160_im <= _T_1159_im;
    _T_1161_re <= _T_1160_re;
    _T_1161_im <= _T_1160_im;
    _T_1162_re <= _T_1161_re;
    _T_1162_im <= _T_1161_im;
    _T_1163_re <= _T_1162_re;
    _T_1163_im <= _T_1162_im;
    _T_1164_re <= _T_1163_re;
    _T_1164_im <= _T_1163_im;
    _T_1165_re <= _T_1164_re;
    _T_1165_im <= _T_1164_im;
    _T_1166_re <= _T_1165_re;
    _T_1166_im <= _T_1165_im;
    _T_1167_re <= _T_1166_re;
    _T_1167_im <= _T_1166_im;
    _T_1168_re <= _T_1167_re;
    _T_1168_im <= _T_1167_im;
    _T_1169_re <= _T_1168_re;
    _T_1169_im <= _T_1168_im;
    _T_1170_re <= _T_1169_re;
    _T_1170_im <= _T_1169_im;
    _T_1171_re <= _T_1170_re;
    _T_1171_im <= _T_1170_im;
    _T_1172_re <= _T_1171_re;
    _T_1172_im <= _T_1171_im;
    _T_1173_re <= _T_1172_re;
    _T_1173_im <= _T_1172_im;
    _T_1174_re <= _T_1173_re;
    _T_1174_im <= _T_1173_im;
    _T_1175_re <= _T_1174_re;
    _T_1175_im <= _T_1174_im;
    _T_1176_re <= _T_1175_re;
    _T_1176_im <= _T_1175_im;
    _T_1177_re <= _T_1176_re;
    _T_1177_im <= _T_1176_im;
    _T_1178_re <= _T_1177_re;
    _T_1178_im <= _T_1177_im;
    _T_1179_re <= _T_1178_re;
    _T_1179_im <= _T_1178_im;
    _T_1180_re <= _T_1179_re;
    _T_1180_im <= _T_1179_im;
    _T_1181_re <= _T_1180_re;
    _T_1181_im <= _T_1180_im;
    _T_1182_re <= _T_1181_re;
    _T_1182_im <= _T_1181_im;
    _T_1183_re <= _T_1182_re;
    _T_1183_im <= _T_1182_im;
    _T_1184_re <= _T_1183_re;
    _T_1184_im <= _T_1183_im;
    _T_1185_re <= _T_1184_re;
    _T_1185_im <= _T_1184_im;
    _T_1186_re <= _T_1185_re;
    _T_1186_im <= _T_1185_im;
    _T_1187_re <= _T_1186_re;
    _T_1187_im <= _T_1186_im;
    _T_1188_re <= _T_1187_re;
    _T_1188_im <= _T_1187_im;
    _T_1189_re <= _T_1188_re;
    _T_1189_im <= _T_1188_im;
    _T_1190_re <= _T_1189_re;
    _T_1190_im <= _T_1189_im;
    _T_1191_re <= _T_1190_re;
    _T_1191_im <= _T_1190_im;
    _T_1192_re <= _T_1191_re;
    _T_1192_im <= _T_1191_im;
    _T_1193_re <= _T_1192_re;
    _T_1193_im <= _T_1192_im;
    _T_1194_re <= _T_1193_re;
    _T_1194_im <= _T_1193_im;
    _T_1195_re <= _T_1194_re;
    _T_1195_im <= _T_1194_im;
    _T_1196_re <= _T_1195_re;
    _T_1196_im <= _T_1195_im;
    _T_1197_re <= _T_1196_re;
    _T_1197_im <= _T_1196_im;
    _T_1198_re <= _T_1197_re;
    _T_1198_im <= _T_1197_im;
    _T_1199_re <= _T_1198_re;
    _T_1199_im <= _T_1198_im;
    _T_1200_re <= _T_1199_re;
    _T_1200_im <= _T_1199_im;
    _T_1201_re <= _T_1200_re;
    _T_1201_im <= _T_1200_im;
    _T_1202_re <= _T_1201_re;
    _T_1202_im <= _T_1201_im;
    _T_1203_re <= _T_1202_re;
    _T_1203_im <= _T_1202_im;
    _T_1204_re <= _T_1203_re;
    _T_1204_im <= _T_1203_im;
    _T_1205_re <= _T_1204_re;
    _T_1205_im <= _T_1204_im;
    _T_1206_re <= _T_1205_re;
    _T_1206_im <= _T_1205_im;
    _T_1207_re <= _T_1206_re;
    _T_1207_im <= _T_1206_im;
    _T_1208_re <= _T_1207_re;
    _T_1208_im <= _T_1207_im;
    _T_1209_re <= _T_1208_re;
    _T_1209_im <= _T_1208_im;
    _T_1210_re <= _T_1209_re;
    _T_1210_im <= _T_1209_im;
    _T_1211_re <= _T_1210_re;
    _T_1211_im <= _T_1210_im;
    _T_1212_re <= _T_1211_re;
    _T_1212_im <= _T_1211_im;
    _T_1213_re <= _T_1212_re;
    _T_1213_im <= _T_1212_im;
    _T_1214_re <= _T_1213_re;
    _T_1214_im <= _T_1213_im;
    _T_1215_re <= _T_1214_re;
    _T_1215_im <= _T_1214_im;
    _T_1216_re <= _T_1215_re;
    _T_1216_im <= _T_1215_im;
    _T_1217_re <= _T_1216_re;
    _T_1217_im <= _T_1216_im;
    _T_1218_re <= _T_1217_re;
    _T_1218_im <= _T_1217_im;
    _T_1219_re <= _T_1218_re;
    _T_1219_im <= _T_1218_im;
    _T_1220_re <= _T_1219_re;
    _T_1220_im <= _T_1219_im;
    _T_1221_re <= _T_1220_re;
    _T_1221_im <= _T_1220_im;
    _T_1222_re <= _T_1221_re;
    _T_1222_im <= _T_1221_im;
    _T_1223_re <= _T_1222_re;
    _T_1223_im <= _T_1222_im;
    _T_1224_re <= _T_1223_re;
    _T_1224_im <= _T_1223_im;
    _T_1225_re <= _T_1224_re;
    _T_1225_im <= _T_1224_im;
    _T_1226_re <= _T_1225_re;
    _T_1226_im <= _T_1225_im;
    _T_1227_re <= _T_1226_re;
    _T_1227_im <= _T_1226_im;
    _T_1228_re <= _T_1227_re;
    _T_1228_im <= _T_1227_im;
    _T_1229_re <= _T_1228_re;
    _T_1229_im <= _T_1228_im;
    _T_1230_re <= _T_1229_re;
    _T_1230_im <= _T_1229_im;
    _T_1231_re <= _T_1230_re;
    _T_1231_im <= _T_1230_im;
    _T_1232_re <= _T_1231_re;
    _T_1232_im <= _T_1231_im;
    _T_1233_re <= _T_1232_re;
    _T_1233_im <= _T_1232_im;
    _T_1234_re <= _T_1233_re;
    _T_1234_im <= _T_1233_im;
    _T_1235_re <= _T_1234_re;
    _T_1235_im <= _T_1234_im;
    _T_1236_re <= _T_1235_re;
    _T_1236_im <= _T_1235_im;
    _T_1237_re <= _T_1236_re;
    _T_1237_im <= _T_1236_im;
    _T_1238_re <= _T_1237_re;
    _T_1238_im <= _T_1237_im;
    _T_1239_re <= _T_1238_re;
    _T_1239_im <= _T_1238_im;
    _T_1240_re <= _T_1239_re;
    _T_1240_im <= _T_1239_im;
    _T_1241_re <= _T_1240_re;
    _T_1241_im <= _T_1240_im;
    _T_1242_re <= _T_1241_re;
    _T_1242_im <= _T_1241_im;
    _T_1243_re <= _T_1242_re;
    _T_1243_im <= _T_1242_im;
    _T_1244_re <= _T_1243_re;
    _T_1244_im <= _T_1243_im;
    _T_1245_re <= _T_1244_re;
    _T_1245_im <= _T_1244_im;
    _T_1246_re <= _T_1245_re;
    _T_1246_im <= _T_1245_im;
    _T_1247_re <= _T_1246_re;
    _T_1247_im <= _T_1246_im;
    _T_1248_re <= _T_1247_re;
    _T_1248_im <= _T_1247_im;
    _T_1249_re <= _T_1248_re;
    _T_1249_im <= _T_1248_im;
    _T_1250_re <= _T_1249_re;
    _T_1250_im <= _T_1249_im;
    _T_1251_re <= _T_1250_re;
    _T_1251_im <= _T_1250_im;
    _T_1252_re <= _T_1251_re;
    _T_1252_im <= _T_1251_im;
    _T_1253_re <= _T_1252_re;
    _T_1253_im <= _T_1252_im;
    _T_1254_re <= _T_1253_re;
    _T_1254_im <= _T_1253_im;
    _T_1255_re <= _T_1254_re;
    _T_1255_im <= _T_1254_im;
    _T_1256_re <= _T_1255_re;
    _T_1256_im <= _T_1255_im;
    _T_1257_re <= _T_1256_re;
    _T_1257_im <= _T_1256_im;
    _T_1258_re <= _T_1257_re;
    _T_1258_im <= _T_1257_im;
    _T_1259_re <= _T_1258_re;
    _T_1259_im <= _T_1258_im;
    _T_1260_re <= _T_1259_re;
    _T_1260_im <= _T_1259_im;
    _T_1261_re <= _T_1260_re;
    _T_1261_im <= _T_1260_im;
    _T_1262_re <= _T_1261_re;
    _T_1262_im <= _T_1261_im;
    _T_1263_re <= _T_1262_re;
    _T_1263_im <= _T_1262_im;
    _T_1264_re <= _T_1263_re;
    _T_1264_im <= _T_1263_im;
    _T_1265_re <= _T_1264_re;
    _T_1265_im <= _T_1264_im;
    _T_1266_re <= _T_1265_re;
    _T_1266_im <= _T_1265_im;
    _T_1267_re <= _T_1266_re;
    _T_1267_im <= _T_1266_im;
    _T_1268_re <= _T_1267_re;
    _T_1268_im <= _T_1267_im;
    _T_1269_re <= _T_1268_re;
    _T_1269_im <= _T_1268_im;
    _T_1270_re <= _T_1269_re;
    _T_1270_im <= _T_1269_im;
    _T_1271_re <= _T_1270_re;
    _T_1271_im <= _T_1270_im;
    _T_1272_re <= _T_1271_re;
    _T_1272_im <= _T_1271_im;
    _T_1273_re <= _T_1272_re;
    _T_1273_im <= _T_1272_im;
    _T_1274_re <= _T_1273_re;
    _T_1274_im <= _T_1273_im;
    _T_1275_re <= _T_1274_re;
    _T_1275_im <= _T_1274_im;
    _T_1276_re <= _T_1275_re;
    _T_1276_im <= _T_1275_im;
    _T_1277_re <= _T_1276_re;
    _T_1277_im <= _T_1276_im;
    _T_1278_re <= _T_1277_re;
    _T_1278_im <= _T_1277_im;
    _T_1279_re <= _T_1278_re;
    _T_1279_im <= _T_1278_im;
    _T_1280_re <= _T_1279_re;
    _T_1280_im <= _T_1279_im;
    _T_1281_re <= _T_1280_re;
    _T_1281_im <= _T_1280_im;
    _T_1282_re <= _T_1281_re;
    _T_1282_im <= _T_1281_im;
    _T_1283_re <= _T_1282_re;
    _T_1283_im <= _T_1282_im;
    _T_1284_re <= _T_1283_re;
    _T_1284_im <= _T_1283_im;
    _T_1285_re <= _T_1284_re;
    _T_1285_im <= _T_1284_im;
    _T_1286_re <= _T_1285_re;
    _T_1286_im <= _T_1285_im;
    _T_1287_re <= _T_1286_re;
    _T_1287_im <= _T_1286_im;
    _T_1288_re <= _T_1287_re;
    _T_1288_im <= _T_1287_im;
    _T_1289_re <= _T_1288_re;
    _T_1289_im <= _T_1288_im;
    _T_1290_re <= _T_1289_re;
    _T_1290_im <= _T_1289_im;
    _T_1291_re <= _T_1290_re;
    _T_1291_im <= _T_1290_im;
    _T_1292_re <= _T_1291_re;
    _T_1292_im <= _T_1291_im;
    _T_1293_re <= _T_1292_re;
    _T_1293_im <= _T_1292_im;
    _T_1294_re <= _T_1293_re;
    _T_1294_im <= _T_1293_im;
    _T_1295_re <= _T_1294_re;
    _T_1295_im <= _T_1294_im;
    _T_1296_re <= _T_1295_re;
    _T_1296_im <= _T_1295_im;
    _T_1297_re <= _T_1296_re;
    _T_1297_im <= _T_1296_im;
    _T_1298_re <= _T_1297_re;
    _T_1298_im <= _T_1297_im;
    _T_1299_re <= _T_1298_re;
    _T_1299_im <= _T_1298_im;
    _T_1300_re <= _T_1299_re;
    _T_1300_im <= _T_1299_im;
    _T_1301_re <= _T_1300_re;
    _T_1301_im <= _T_1300_im;
    _T_1302_re <= _T_1301_re;
    _T_1302_im <= _T_1301_im;
    _T_1303_re <= _T_1302_re;
    _T_1303_im <= _T_1302_im;
    _T_1304_re <= _T_1303_re;
    _T_1304_im <= _T_1303_im;
    _T_1305_re <= _T_1304_re;
    _T_1305_im <= _T_1304_im;
    _T_1306_re <= _T_1305_re;
    _T_1306_im <= _T_1305_im;
    _T_1307_re <= _T_1306_re;
    _T_1307_im <= _T_1306_im;
    _T_1308_re <= _T_1307_re;
    _T_1308_im <= _T_1307_im;
    _T_1309_re <= _T_1308_re;
    _T_1309_im <= _T_1308_im;
    _T_1310_re <= _T_1309_re;
    _T_1310_im <= _T_1309_im;
    _T_1311_re <= _T_1310_re;
    _T_1311_im <= _T_1310_im;
    _T_1312_re <= _T_1311_re;
    _T_1312_im <= _T_1311_im;
    _T_1313_re <= _T_1312_re;
    _T_1313_im <= _T_1312_im;
    _T_1314_re <= _T_1313_re;
    _T_1314_im <= _T_1313_im;
    _T_1315_re <= _T_1314_re;
    _T_1315_im <= _T_1314_im;
    _T_1316_re <= _T_1315_re;
    _T_1316_im <= _T_1315_im;
    _T_1317_re <= _T_1316_re;
    _T_1317_im <= _T_1316_im;
    _T_1318_re <= _T_1317_re;
    _T_1318_im <= _T_1317_im;
    _T_1319_re <= _T_1318_re;
    _T_1319_im <= _T_1318_im;
    _T_1320_re <= _T_1319_re;
    _T_1320_im <= _T_1319_im;
    _T_1321_re <= _T_1320_re;
    _T_1321_im <= _T_1320_im;
    _T_1322_re <= _T_1321_re;
    _T_1322_im <= _T_1321_im;
    _T_1323_re <= _T_1322_re;
    _T_1323_im <= _T_1322_im;
    _T_1324_re <= _T_1323_re;
    _T_1324_im <= _T_1323_im;
    _T_1325_re <= _T_1324_re;
    _T_1325_im <= _T_1324_im;
    _T_1326_re <= _T_1325_re;
    _T_1326_im <= _T_1325_im;
    _T_1327_re <= _T_1326_re;
    _T_1327_im <= _T_1326_im;
    _T_1328_re <= _T_1327_re;
    _T_1328_im <= _T_1327_im;
    _T_1329_re <= _T_1328_re;
    _T_1329_im <= _T_1328_im;
    _T_1330_re <= _T_1329_re;
    _T_1330_im <= _T_1329_im;
    _T_1331_re <= _T_1330_re;
    _T_1331_im <= _T_1330_im;
    _T_1332_re <= _T_1331_re;
    _T_1332_im <= _T_1331_im;
    _T_1333_re <= _T_1332_re;
    _T_1333_im <= _T_1332_im;
    _T_1334_re <= _T_1333_re;
    _T_1334_im <= _T_1333_im;
    _T_1335_re <= _T_1334_re;
    _T_1335_im <= _T_1334_im;
    _T_1336_re <= _T_1335_re;
    _T_1336_im <= _T_1335_im;
    _T_1337_re <= _T_1336_re;
    _T_1337_im <= _T_1336_im;
    _T_1338_re <= _T_1337_re;
    _T_1338_im <= _T_1337_im;
    _T_1339_re <= _T_1338_re;
    _T_1339_im <= _T_1338_im;
    _T_1340_re <= _T_1339_re;
    _T_1340_im <= _T_1339_im;
    _T_1341_re <= _T_1340_re;
    _T_1341_im <= _T_1340_im;
    _T_1342_re <= _T_1341_re;
    _T_1342_im <= _T_1341_im;
    _T_1343_re <= _T_1342_re;
    _T_1343_im <= _T_1342_im;
    _T_1344_re <= _T_1343_re;
    _T_1344_im <= _T_1343_im;
    _T_1345_re <= _T_1344_re;
    _T_1345_im <= _T_1344_im;
    _T_1346_re <= _T_1345_re;
    _T_1346_im <= _T_1345_im;
    _T_1347_re <= _T_1346_re;
    _T_1347_im <= _T_1346_im;
    _T_1348_re <= _T_1347_re;
    _T_1348_im <= _T_1347_im;
    _T_1349_re <= _T_1348_re;
    _T_1349_im <= _T_1348_im;
    _T_1350_re <= _T_1349_re;
    _T_1350_im <= _T_1349_im;
    _T_1351_re <= _T_1350_re;
    _T_1351_im <= _T_1350_im;
    _T_1352_re <= _T_1351_re;
    _T_1352_im <= _T_1351_im;
    _T_1353_re <= _T_1352_re;
    _T_1353_im <= _T_1352_im;
    _T_1354_re <= _T_1353_re;
    _T_1354_im <= _T_1353_im;
    _T_1355_re <= _T_1354_re;
    _T_1355_im <= _T_1354_im;
    _T_1356_re <= _T_1355_re;
    _T_1356_im <= _T_1355_im;
    _T_1357_re <= _T_1356_re;
    _T_1357_im <= _T_1356_im;
    _T_1358_re <= _T_1357_re;
    _T_1358_im <= _T_1357_im;
    _T_1359_re <= _T_1358_re;
    _T_1359_im <= _T_1358_im;
    _T_1360_re <= _T_1359_re;
    _T_1360_im <= _T_1359_im;
    _T_1361_re <= _T_1360_re;
    _T_1361_im <= _T_1360_im;
    _T_1362_re <= _T_1361_re;
    _T_1362_im <= _T_1361_im;
    _T_1363_re <= _T_1362_re;
    _T_1363_im <= _T_1362_im;
    _T_1364_re <= _T_1363_re;
    _T_1364_im <= _T_1363_im;
    _T_1365_re <= _T_1364_re;
    _T_1365_im <= _T_1364_im;
    _T_1366_re <= _T_1365_re;
    _T_1366_im <= _T_1365_im;
    _T_1367_re <= _T_1366_re;
    _T_1367_im <= _T_1366_im;
    _T_1368_re <= _T_1367_re;
    _T_1368_im <= _T_1367_im;
    _T_1369_re <= _T_1368_re;
    _T_1369_im <= _T_1368_im;
    _T_1370_re <= _T_1369_re;
    _T_1370_im <= _T_1369_im;
    _T_1371_re <= _T_1370_re;
    _T_1371_im <= _T_1370_im;
    _T_1372_re <= _T_1371_re;
    _T_1372_im <= _T_1371_im;
    _T_1373_re <= _T_1372_re;
    _T_1373_im <= _T_1372_im;
    _T_1374_re <= _T_1373_re;
    _T_1374_im <= _T_1373_im;
    _T_1375_re <= _T_1374_re;
    _T_1375_im <= _T_1374_im;
    _T_1376_re <= _T_1375_re;
    _T_1376_im <= _T_1375_im;
    _T_1377_re <= _T_1376_re;
    _T_1377_im <= _T_1376_im;
    _T_1378_re <= _T_1377_re;
    _T_1378_im <= _T_1377_im;
    _T_1379_re <= _T_1378_re;
    _T_1379_im <= _T_1378_im;
    _T_1380_re <= _T_1379_re;
    _T_1380_im <= _T_1379_im;
    _T_1381_re <= _T_1380_re;
    _T_1381_im <= _T_1380_im;
    _T_1382_re <= _T_1381_re;
    _T_1382_im <= _T_1381_im;
    _T_1383_re <= _T_1382_re;
    _T_1383_im <= _T_1382_im;
    _T_1384_re <= _T_1383_re;
    _T_1384_im <= _T_1383_im;
    _T_1385_re <= _T_1384_re;
    _T_1385_im <= _T_1384_im;
    _T_1386_re <= _T_1385_re;
    _T_1386_im <= _T_1385_im;
    _T_1387_re <= _T_1386_re;
    _T_1387_im <= _T_1386_im;
    _T_1388_re <= _T_1387_re;
    _T_1388_im <= _T_1387_im;
    _T_1389_re <= _T_1388_re;
    _T_1389_im <= _T_1388_im;
    _T_1390_re <= _T_1389_re;
    _T_1390_im <= _T_1389_im;
    _T_1391_re <= _T_1390_re;
    _T_1391_im <= _T_1390_im;
    _T_1392_re <= _T_1391_re;
    _T_1392_im <= _T_1391_im;
    _T_1393_re <= _T_1392_re;
    _T_1393_im <= _T_1392_im;
    _T_1394_re <= _T_1393_re;
    _T_1394_im <= _T_1393_im;
    _T_1395_re <= _T_1394_re;
    _T_1395_im <= _T_1394_im;
    _T_1396_re <= _T_1395_re;
    _T_1396_im <= _T_1395_im;
    _T_1397_re <= _T_1396_re;
    _T_1397_im <= _T_1396_im;
    _T_1398_re <= _T_1397_re;
    _T_1398_im <= _T_1397_im;
    _T_1399_re <= _T_1398_re;
    _T_1399_im <= _T_1398_im;
    _T_1400_re <= _T_1399_re;
    _T_1400_im <= _T_1399_im;
    _T_1401_re <= _T_1400_re;
    _T_1401_im <= _T_1400_im;
    _T_1402_re <= _T_1401_re;
    _T_1402_im <= _T_1401_im;
    _T_1403_re <= _T_1402_re;
    _T_1403_im <= _T_1402_im;
    _T_1404_re <= _T_1403_re;
    _T_1404_im <= _T_1403_im;
    _T_1405_re <= _T_1404_re;
    _T_1405_im <= _T_1404_im;
    _T_1406_re <= _T_1405_re;
    _T_1406_im <= _T_1405_im;
    _T_1407_re <= _T_1406_re;
    _T_1407_im <= _T_1406_im;
    _T_1408_re <= _T_1407_re;
    _T_1408_im <= _T_1407_im;
    _T_1409_re <= _T_1408_re;
    _T_1409_im <= _T_1408_im;
    _T_1410_re <= _T_1409_re;
    _T_1410_im <= _T_1409_im;
    _T_1411_re <= _T_1410_re;
    _T_1411_im <= _T_1410_im;
    _T_1412_re <= _T_1411_re;
    _T_1412_im <= _T_1411_im;
    _T_1413_re <= _T_1412_re;
    _T_1413_im <= _T_1412_im;
    _T_1414_re <= _T_1413_re;
    _T_1414_im <= _T_1413_im;
    _T_1415_re <= _T_1414_re;
    _T_1415_im <= _T_1414_im;
    _T_1416_re <= _T_1415_re;
    _T_1416_im <= _T_1415_im;
    _T_1417_re <= _T_1416_re;
    _T_1417_im <= _T_1416_im;
    _T_1418_re <= _T_1417_re;
    _T_1418_im <= _T_1417_im;
    _T_1419_re <= _T_1418_re;
    _T_1419_im <= _T_1418_im;
    _T_1420_re <= _T_1419_re;
    _T_1420_im <= _T_1419_im;
    _T_1421_re <= _T_1420_re;
    _T_1421_im <= _T_1420_im;
    _T_1422_re <= _T_1421_re;
    _T_1422_im <= _T_1421_im;
    _T_1423_re <= _T_1422_re;
    _T_1423_im <= _T_1422_im;
    _T_1424_re <= _T_1423_re;
    _T_1424_im <= _T_1423_im;
    _T_1425_re <= _T_1424_re;
    _T_1425_im <= _T_1424_im;
    _T_1426_re <= _T_1425_re;
    _T_1426_im <= _T_1425_im;
    _T_1427_re <= _T_1426_re;
    _T_1427_im <= _T_1426_im;
    _T_1428_re <= _T_1427_re;
    _T_1428_im <= _T_1427_im;
    _T_1429_re <= _T_1428_re;
    _T_1429_im <= _T_1428_im;
    _T_1430_re <= _T_1429_re;
    _T_1430_im <= _T_1429_im;
    _T_1431_re <= _T_1430_re;
    _T_1431_im <= _T_1430_im;
    _T_1432_re <= _T_1431_re;
    _T_1432_im <= _T_1431_im;
    _T_1433_re <= _T_1432_re;
    _T_1433_im <= _T_1432_im;
    _T_1434_re <= _T_1433_re;
    _T_1434_im <= _T_1433_im;
    _T_1435_re <= _T_1434_re;
    _T_1435_im <= _T_1434_im;
    _T_1436_re <= _T_1435_re;
    _T_1436_im <= _T_1435_im;
    _T_1437_re <= _T_1436_re;
    _T_1437_im <= _T_1436_im;
    _T_1438_re <= _T_1437_re;
    _T_1438_im <= _T_1437_im;
    _T_1439_re <= _T_1438_re;
    _T_1439_im <= _T_1438_im;
    _T_1440_re <= _T_1439_re;
    _T_1440_im <= _T_1439_im;
    _T_1441_re <= _T_1440_re;
    _T_1441_im <= _T_1440_im;
    _T_1442_re <= _T_1441_re;
    _T_1442_im <= _T_1441_im;
    _T_1443_re <= _T_1442_re;
    _T_1443_im <= _T_1442_im;
    _T_1444_re <= _T_1443_re;
    _T_1444_im <= _T_1443_im;
    _T_1445_re <= _T_1444_re;
    _T_1445_im <= _T_1444_im;
    _T_1446_re <= _T_1445_re;
    _T_1446_im <= _T_1445_im;
    _T_1447_re <= _T_1446_re;
    _T_1447_im <= _T_1446_im;
    _T_1448_re <= _T_1447_re;
    _T_1448_im <= _T_1447_im;
    _T_1449_re <= _T_1448_re;
    _T_1449_im <= _T_1448_im;
    _T_1450_re <= _T_1449_re;
    _T_1450_im <= _T_1449_im;
    _T_1451_re <= _T_1450_re;
    _T_1451_im <= _T_1450_im;
    _T_1452_re <= _T_1451_re;
    _T_1452_im <= _T_1451_im;
    _T_1453_re <= _T_1452_re;
    _T_1453_im <= _T_1452_im;
    _T_1454_re <= _T_1453_re;
    _T_1454_im <= _T_1453_im;
    _T_1455_re <= _T_1454_re;
    _T_1455_im <= _T_1454_im;
    _T_1456_re <= _T_1455_re;
    _T_1456_im <= _T_1455_im;
    _T_1457_re <= _T_1456_re;
    _T_1457_im <= _T_1456_im;
    _T_1458_re <= _T_1457_re;
    _T_1458_im <= _T_1457_im;
    _T_1459_re <= _T_1458_re;
    _T_1459_im <= _T_1458_im;
    _T_1460_re <= _T_1459_re;
    _T_1460_im <= _T_1459_im;
    _T_1461_re <= _T_1460_re;
    _T_1461_im <= _T_1460_im;
    _T_1462_re <= _T_1461_re;
    _T_1462_im <= _T_1461_im;
    _T_1463_re <= _T_1462_re;
    _T_1463_im <= _T_1462_im;
    _T_1464_re <= _T_1463_re;
    _T_1464_im <= _T_1463_im;
    _T_1465_re <= _T_1464_re;
    _T_1465_im <= _T_1464_im;
    _T_1466_re <= _T_1465_re;
    _T_1466_im <= _T_1465_im;
    _T_1467_re <= _T_1466_re;
    _T_1467_im <= _T_1466_im;
    _T_1468_re <= _T_1467_re;
    _T_1468_im <= _T_1467_im;
    _T_1469_re <= _T_1468_re;
    _T_1469_im <= _T_1468_im;
    _T_1470_re <= _T_1469_re;
    _T_1470_im <= _T_1469_im;
    _T_1471_re <= _T_1470_re;
    _T_1471_im <= _T_1470_im;
    _T_1472_re <= _T_1471_re;
    _T_1472_im <= _T_1471_im;
    _T_1473_re <= _T_1472_re;
    _T_1473_im <= _T_1472_im;
    _T_1474_re <= _T_1473_re;
    _T_1474_im <= _T_1473_im;
    _T_1475_re <= _T_1474_re;
    _T_1475_im <= _T_1474_im;
    _T_1476_re <= _T_1475_re;
    _T_1476_im <= _T_1475_im;
    _T_1477_re <= _T_1476_re;
    _T_1477_im <= _T_1476_im;
    _T_1478_re <= _T_1477_re;
    _T_1478_im <= _T_1477_im;
    _T_1479_re <= _T_1478_re;
    _T_1479_im <= _T_1478_im;
    _T_1480_re <= _T_1479_re;
    _T_1480_im <= _T_1479_im;
    _T_1481_re <= _T_1480_re;
    _T_1481_im <= _T_1480_im;
    _T_1482_re <= _T_1481_re;
    _T_1482_im <= _T_1481_im;
    _T_1483_re <= _T_1482_re;
    _T_1483_im <= _T_1482_im;
    _T_1484_re <= _T_1483_re;
    _T_1484_im <= _T_1483_im;
    _T_1485_re <= _T_1484_re;
    _T_1485_im <= _T_1484_im;
    _T_1486_re <= _T_1485_re;
    _T_1486_im <= _T_1485_im;
    _T_1487_re <= _T_1486_re;
    _T_1487_im <= _T_1486_im;
    _T_1488_re <= _T_1487_re;
    _T_1488_im <= _T_1487_im;
    _T_1489_re <= _T_1488_re;
    _T_1489_im <= _T_1488_im;
    _T_1490_re <= _T_1489_re;
    _T_1490_im <= _T_1489_im;
    _T_1491_re <= _T_1490_re;
    _T_1491_im <= _T_1490_im;
    _T_1492_re <= _T_1491_re;
    _T_1492_im <= _T_1491_im;
    _T_1493_re <= _T_1492_re;
    _T_1493_im <= _T_1492_im;
    _T_1494_re <= _T_1493_re;
    _T_1494_im <= _T_1493_im;
    _T_1495_re <= _T_1494_re;
    _T_1495_im <= _T_1494_im;
    _T_1496_re <= _T_1495_re;
    _T_1496_im <= _T_1495_im;
    _T_1497_re <= _T_1496_re;
    _T_1497_im <= _T_1496_im;
    _T_1498_re <= _T_1497_re;
    _T_1498_im <= _T_1497_im;
    _T_1499_re <= _T_1498_re;
    _T_1499_im <= _T_1498_im;
    _T_1500_re <= _T_1499_re;
    _T_1500_im <= _T_1499_im;
    _T_1501_re <= _T_1500_re;
    _T_1501_im <= _T_1500_im;
    _T_1502_re <= _T_1501_re;
    _T_1502_im <= _T_1501_im;
    _T_1503_re <= _T_1502_re;
    _T_1503_im <= _T_1502_im;
    _T_1504_re <= _T_1503_re;
    _T_1504_im <= _T_1503_im;
    _T_1505_re <= _T_1504_re;
    _T_1505_im <= _T_1504_im;
    _T_1506_re <= _T_1505_re;
    _T_1506_im <= _T_1505_im;
    _T_1507_re <= _T_1506_re;
    _T_1507_im <= _T_1506_im;
    _T_1508_re <= _T_1507_re;
    _T_1508_im <= _T_1507_im;
    _T_1509_re <= _T_1508_re;
    _T_1509_im <= _T_1508_im;
    _T_1510_re <= _T_1509_re;
    _T_1510_im <= _T_1509_im;
    _T_1511_re <= _T_1510_re;
    _T_1511_im <= _T_1510_im;
    _T_1512_re <= _T_1511_re;
    _T_1512_im <= _T_1511_im;
    _T_1513_re <= _T_1512_re;
    _T_1513_im <= _T_1512_im;
    _T_1514_re <= _T_1513_re;
    _T_1514_im <= _T_1513_im;
    _T_1515_re <= _T_1514_re;
    _T_1515_im <= _T_1514_im;
    _T_1516_re <= _T_1515_re;
    _T_1516_im <= _T_1515_im;
    _T_1517_re <= _T_1516_re;
    _T_1517_im <= _T_1516_im;
    _T_1518_re <= _T_1517_re;
    _T_1518_im <= _T_1517_im;
    _T_1519_re <= _T_1518_re;
    _T_1519_im <= _T_1518_im;
    _T_1520_re <= _T_1519_re;
    _T_1520_im <= _T_1519_im;
    _T_1521_re <= _T_1520_re;
    _T_1521_im <= _T_1520_im;
    _T_1522_re <= _T_1521_re;
    _T_1522_im <= _T_1521_im;
    _T_1523_re <= _T_1522_re;
    _T_1523_im <= _T_1522_im;
    _T_1524_re <= _T_1523_re;
    _T_1524_im <= _T_1523_im;
    _T_1525_re <= _T_1524_re;
    _T_1525_im <= _T_1524_im;
    _T_1526_re <= _T_1525_re;
    _T_1526_im <= _T_1525_im;
    _T_1527_re <= _T_1526_re;
    _T_1527_im <= _T_1526_im;
    _T_1528_re <= _T_1527_re;
    _T_1528_im <= _T_1527_im;
    _T_1529_re <= _T_1528_re;
    _T_1529_im <= _T_1528_im;
    _T_1530_re <= _T_1529_re;
    _T_1530_im <= _T_1529_im;
    _T_1531_re <= _T_1530_re;
    _T_1531_im <= _T_1530_im;
    _T_1532_re <= _T_1531_re;
    _T_1532_im <= _T_1531_im;
    _T_1533_re <= _T_1532_re;
    _T_1533_im <= _T_1532_im;
    _T_1534_re <= _T_1533_re;
    _T_1534_im <= _T_1533_im;
    _T_1535_re <= _T_1534_re;
    _T_1535_im <= _T_1534_im;
    _T_1536_re <= _T_1535_re;
    _T_1536_im <= _T_1535_im;
    _T_1537_re <= _T_1536_re;
    _T_1537_im <= _T_1536_im;
    _T_1538_re <= _T_1537_re;
    _T_1538_im <= _T_1537_im;
    _T_1539_re <= _T_1538_re;
    _T_1539_im <= _T_1538_im;
    _T_1540_re <= _T_1539_re;
    _T_1540_im <= _T_1539_im;
    _T_1541_re <= _T_1540_re;
    _T_1541_im <= _T_1540_im;
    _T_1542_re <= _T_1541_re;
    _T_1542_im <= _T_1541_im;
    _T_1543_re <= _T_1542_re;
    _T_1543_im <= _T_1542_im;
    _T_1544_re <= _T_1543_re;
    _T_1544_im <= _T_1543_im;
    _T_1545_re <= _T_1544_re;
    _T_1545_im <= _T_1544_im;
    _T_1546_re <= _T_1545_re;
    _T_1546_im <= _T_1545_im;
    _T_1547_re <= _T_1546_re;
    _T_1547_im <= _T_1546_im;
    _T_1548_re <= _T_1547_re;
    _T_1548_im <= _T_1547_im;
    _T_1549_re <= _T_1548_re;
    _T_1549_im <= _T_1548_im;
    _T_1550_re <= _T_1549_re;
    _T_1550_im <= _T_1549_im;
    _T_1551_re <= _T_1550_re;
    _T_1551_im <= _T_1550_im;
    _T_1552_re <= _T_1551_re;
    _T_1552_im <= _T_1551_im;
    _T_1553_re <= _T_1552_re;
    _T_1553_im <= _T_1552_im;
    _T_1554_re <= _T_1553_re;
    _T_1554_im <= _T_1553_im;
    _T_1555_re <= _T_1554_re;
    _T_1555_im <= _T_1554_im;
    _T_1556_re <= _T_1555_re;
    _T_1556_im <= _T_1555_im;
    _T_1557_re <= _T_1556_re;
    _T_1557_im <= _T_1556_im;
    _T_1558_re <= _T_1557_re;
    _T_1558_im <= _T_1557_im;
    _T_1559_re <= _T_1558_re;
    _T_1559_im <= _T_1558_im;
    _T_1560_re <= _T_1559_re;
    _T_1560_im <= _T_1559_im;
    _T_1561_re <= _T_1560_re;
    _T_1561_im <= _T_1560_im;
    _T_1562_re <= _T_1561_re;
    _T_1562_im <= _T_1561_im;
    _T_1563_re <= _T_1562_re;
    _T_1563_im <= _T_1562_im;
    _T_1564_re <= _T_1563_re;
    _T_1564_im <= _T_1563_im;
    _T_1565_re <= _T_1564_re;
    _T_1565_im <= _T_1564_im;
    _T_1566_re <= _T_1565_re;
    _T_1566_im <= _T_1565_im;
    _T_1567_re <= _T_1566_re;
    _T_1567_im <= _T_1566_im;
    _T_1568_re <= _T_1567_re;
    _T_1568_im <= _T_1567_im;
    _T_1569_re <= _T_1568_re;
    _T_1569_im <= _T_1568_im;
    _T_1570_re <= _T_1569_re;
    _T_1570_im <= _T_1569_im;
    _T_1571_re <= _T_1570_re;
    _T_1571_im <= _T_1570_im;
    _T_1572_re <= _T_1571_re;
    _T_1572_im <= _T_1571_im;
    _T_1573_re <= _T_1572_re;
    _T_1573_im <= _T_1572_im;
    _T_1574_re <= _T_1573_re;
    _T_1574_im <= _T_1573_im;
    _T_1575_re <= _T_1574_re;
    _T_1575_im <= _T_1574_im;
    _T_1576_re <= _T_1575_re;
    _T_1576_im <= _T_1575_im;
    _T_1577_re <= _T_1576_re;
    _T_1577_im <= _T_1576_im;
    _T_1578_re <= _T_1577_re;
    _T_1578_im <= _T_1577_im;
    _T_1579_re <= _T_1578_re;
    _T_1579_im <= _T_1578_im;
    _T_1580_re <= _T_1579_re;
    _T_1580_im <= _T_1579_im;
    _T_1581_re <= _T_1580_re;
    _T_1581_im <= _T_1580_im;
    _T_1582_re <= _T_1581_re;
    _T_1582_im <= _T_1581_im;
    _T_1583_re <= _T_1582_re;
    _T_1583_im <= _T_1582_im;
    _T_1584_re <= _T_1583_re;
    _T_1584_im <= _T_1583_im;
    _T_1585_re <= _T_1584_re;
    _T_1585_im <= _T_1584_im;
    _T_1586_re <= _T_1585_re;
    _T_1586_im <= _T_1585_im;
    _T_1587_re <= _T_1586_re;
    _T_1587_im <= _T_1586_im;
    _T_1588_re <= _T_1587_re;
    _T_1588_im <= _T_1587_im;
    _T_1589_re <= _T_1588_re;
    _T_1589_im <= _T_1588_im;
    _T_1590_re <= _T_1589_re;
    _T_1590_im <= _T_1589_im;
    _T_1591_re <= _T_1590_re;
    _T_1591_im <= _T_1590_im;
    _T_1592_re <= _T_1591_re;
    _T_1592_im <= _T_1591_im;
    _T_1593_re <= _T_1592_re;
    _T_1593_im <= _T_1592_im;
    _T_1594_re <= _T_1593_re;
    _T_1594_im <= _T_1593_im;
    _T_1595_re <= _T_1594_re;
    _T_1595_im <= _T_1594_im;
    _T_1596_re <= _T_1595_re;
    _T_1596_im <= _T_1595_im;
    _T_1597_re <= _T_1596_re;
    _T_1597_im <= _T_1596_im;
    _T_1598_re <= _T_1597_re;
    _T_1598_im <= _T_1597_im;
    _T_1599_re <= _T_1598_re;
    _T_1599_im <= _T_1598_im;
    _T_1600_re <= _T_1599_re;
    _T_1600_im <= _T_1599_im;
    _T_1601_re <= _T_1600_re;
    _T_1601_im <= _T_1600_im;
    _T_1602_re <= _T_1601_re;
    _T_1602_im <= _T_1601_im;
    _T_1603_re <= _T_1602_re;
    _T_1603_im <= _T_1602_im;
    _T_1604_re <= _T_1603_re;
    _T_1604_im <= _T_1603_im;
    _T_1605_re <= _T_1604_re;
    _T_1605_im <= _T_1604_im;
    _T_1606_re <= _T_1605_re;
    _T_1606_im <= _T_1605_im;
    _T_1607_re <= _T_1606_re;
    _T_1607_im <= _T_1606_im;
    _T_1608_re <= _T_1607_re;
    _T_1608_im <= _T_1607_im;
    _T_1609_re <= _T_1608_re;
    _T_1609_im <= _T_1608_im;
    _T_1610_re <= _T_1609_re;
    _T_1610_im <= _T_1609_im;
    _T_1611_re <= _T_1610_re;
    _T_1611_im <= _T_1610_im;
    _T_1612_re <= _T_1611_re;
    _T_1612_im <= _T_1611_im;
    _T_1613_re <= _T_1612_re;
    _T_1613_im <= _T_1612_im;
    _T_1614_re <= _T_1613_re;
    _T_1614_im <= _T_1613_im;
    _T_1615_re <= _T_1614_re;
    _T_1615_im <= _T_1614_im;
    _T_1616_re <= _T_1615_re;
    _T_1616_im <= _T_1615_im;
    _T_1617_re <= _T_1616_re;
    _T_1617_im <= _T_1616_im;
    _T_1618_re <= _T_1617_re;
    _T_1618_im <= _T_1617_im;
    _T_1619_re <= _T_1618_re;
    _T_1619_im <= _T_1618_im;
    _T_1620_re <= _T_1619_re;
    _T_1620_im <= _T_1619_im;
    _T_1621_re <= _T_1620_re;
    _T_1621_im <= _T_1620_im;
    _T_1622_re <= _T_1621_re;
    _T_1622_im <= _T_1621_im;
    _T_1623_re <= _T_1622_re;
    _T_1623_im <= _T_1622_im;
    _T_1624_re <= _T_1623_re;
    _T_1624_im <= _T_1623_im;
    _T_1625_re <= _T_1624_re;
    _T_1625_im <= _T_1624_im;
    _T_1626_re <= _T_1625_re;
    _T_1626_im <= _T_1625_im;
    _T_1627_re <= _T_1626_re;
    _T_1627_im <= _T_1626_im;
    _T_1628_re <= _T_1627_re;
    _T_1628_im <= _T_1627_im;
    _T_1629_re <= _T_1628_re;
    _T_1629_im <= _T_1628_im;
    _T_1630_re <= _T_1629_re;
    _T_1630_im <= _T_1629_im;
    _T_1631_re <= _T_1630_re;
    _T_1631_im <= _T_1630_im;
    _T_1632_re <= _T_1631_re;
    _T_1632_im <= _T_1631_im;
    _T_1633_re <= _T_1632_re;
    _T_1633_im <= _T_1632_im;
    _T_1634_re <= _T_1633_re;
    _T_1634_im <= _T_1633_im;
    _T_1635_re <= _T_1634_re;
    _T_1635_im <= _T_1634_im;
    _T_1636_re <= _T_1635_re;
    _T_1636_im <= _T_1635_im;
    _T_1637_re <= _T_1636_re;
    _T_1637_im <= _T_1636_im;
    _T_1638_re <= _T_1637_re;
    _T_1638_im <= _T_1637_im;
    _T_1639_re <= _T_1638_re;
    _T_1639_im <= _T_1638_im;
    _T_1640_re <= _T_1639_re;
    _T_1640_im <= _T_1639_im;
    _T_1641_re <= _T_1640_re;
    _T_1641_im <= _T_1640_im;
    _T_1642_re <= _T_1641_re;
    _T_1642_im <= _T_1641_im;
    _T_1643_re <= _T_1642_re;
    _T_1643_im <= _T_1642_im;
    _T_1644_re <= _T_1643_re;
    _T_1644_im <= _T_1643_im;
    _T_1645_re <= _T_1644_re;
    _T_1645_im <= _T_1644_im;
    _T_1646_re <= _T_1645_re;
    _T_1646_im <= _T_1645_im;
    _T_1647_re <= _T_1646_re;
    _T_1647_im <= _T_1646_im;
    _T_1648_re <= _T_1647_re;
    _T_1648_im <= _T_1647_im;
    _T_1649_re <= _T_1648_re;
    _T_1649_im <= _T_1648_im;
    _T_1650_re <= _T_1649_re;
    _T_1650_im <= _T_1649_im;
    _T_1651_re <= _T_1650_re;
    _T_1651_im <= _T_1650_im;
    _T_1652_re <= _T_1651_re;
    _T_1652_im <= _T_1651_im;
    _T_1653_re <= _T_1652_re;
    _T_1653_im <= _T_1652_im;
    _T_1654_re <= _T_1653_re;
    _T_1654_im <= _T_1653_im;
    _T_1655_re <= _T_1654_re;
    _T_1655_im <= _T_1654_im;
    _T_1656_re <= _T_1655_re;
    _T_1656_im <= _T_1655_im;
    _T_1657_re <= _T_1656_re;
    _T_1657_im <= _T_1656_im;
    _T_1658_re <= _T_1657_re;
    _T_1658_im <= _T_1657_im;
    _T_1659_re <= _T_1658_re;
    _T_1659_im <= _T_1658_im;
    _T_1660_re <= _T_1659_re;
    _T_1660_im <= _T_1659_im;
    _T_1661_re <= _T_1660_re;
    _T_1661_im <= _T_1660_im;
    _T_1662_re <= _T_1661_re;
    _T_1662_im <= _T_1661_im;
    _T_1663_re <= _T_1662_re;
    _T_1663_im <= _T_1662_im;
    _T_1664_re <= _T_1663_re;
    _T_1664_im <= _T_1663_im;
    _T_1665_re <= _T_1664_re;
    _T_1665_im <= _T_1664_im;
    _T_1666_re <= _T_1665_re;
    _T_1666_im <= _T_1665_im;
    _T_1667_re <= _T_1666_re;
    _T_1667_im <= _T_1666_im;
    _T_1668_re <= _T_1667_re;
    _T_1668_im <= _T_1667_im;
    _T_1669_re <= _T_1668_re;
    _T_1669_im <= _T_1668_im;
    _T_1670_re <= _T_1669_re;
    _T_1670_im <= _T_1669_im;
    _T_1671_re <= _T_1670_re;
    _T_1671_im <= _T_1670_im;
    _T_1672_re <= _T_1671_re;
    _T_1672_im <= _T_1671_im;
    _T_1673_re <= _T_1672_re;
    _T_1673_im <= _T_1672_im;
    _T_1674_re <= _T_1673_re;
    _T_1674_im <= _T_1673_im;
    _T_1675_re <= _T_1674_re;
    _T_1675_im <= _T_1674_im;
    _T_1676_re <= _T_1675_re;
    _T_1676_im <= _T_1675_im;
    _T_1677_re <= _T_1676_re;
    _T_1677_im <= _T_1676_im;
    _T_1678_re <= _T_1677_re;
    _T_1678_im <= _T_1677_im;
    _T_1679_re <= _T_1678_re;
    _T_1679_im <= _T_1678_im;
    _T_1680_re <= _T_1679_re;
    _T_1680_im <= _T_1679_im;
    _T_1681_re <= _T_1680_re;
    _T_1681_im <= _T_1680_im;
    _T_1682_re <= _T_1681_re;
    _T_1682_im <= _T_1681_im;
    _T_1683_re <= _T_1682_re;
    _T_1683_im <= _T_1682_im;
    _T_1684_re <= _T_1683_re;
    _T_1684_im <= _T_1683_im;
    _T_1685_re <= _T_1684_re;
    _T_1685_im <= _T_1684_im;
    _T_1686_re <= _T_1685_re;
    _T_1686_im <= _T_1685_im;
    _T_1687_re <= _T_1686_re;
    _T_1687_im <= _T_1686_im;
    _T_1688_re <= _T_1687_re;
    _T_1688_im <= _T_1687_im;
    _T_1689_re <= _T_1688_re;
    _T_1689_im <= _T_1688_im;
    _T_1690_re <= _T_1689_re;
    _T_1690_im <= _T_1689_im;
    _T_1691_re <= _T_1690_re;
    _T_1691_im <= _T_1690_im;
    _T_1692_re <= _T_1691_re;
    _T_1692_im <= _T_1691_im;
    _T_1693_re <= _T_1692_re;
    _T_1693_im <= _T_1692_im;
    _T_1694_re <= _T_1693_re;
    _T_1694_im <= _T_1693_im;
    _T_1695_re <= _T_1694_re;
    _T_1695_im <= _T_1694_im;
    _T_1696_re <= _T_1695_re;
    _T_1696_im <= _T_1695_im;
    _T_1697_re <= _T_1696_re;
    _T_1697_im <= _T_1696_im;
    _T_1698_re <= _T_1697_re;
    _T_1698_im <= _T_1697_im;
    _T_1699_re <= _T_1698_re;
    _T_1699_im <= _T_1698_im;
    _T_1700_re <= _T_1699_re;
    _T_1700_im <= _T_1699_im;
    _T_1701_re <= _T_1700_re;
    _T_1701_im <= _T_1700_im;
    _T_1702_re <= _T_1701_re;
    _T_1702_im <= _T_1701_im;
    _T_1703_re <= _T_1702_re;
    _T_1703_im <= _T_1702_im;
    _T_1704_re <= _T_1703_re;
    _T_1704_im <= _T_1703_im;
    _T_1705_re <= _T_1704_re;
    _T_1705_im <= _T_1704_im;
    _T_1706_re <= _T_1705_re;
    _T_1706_im <= _T_1705_im;
    _T_1707_re <= _T_1706_re;
    _T_1707_im <= _T_1706_im;
    _T_1708_re <= _T_1707_re;
    _T_1708_im <= _T_1707_im;
    _T_1709_re <= _T_1708_re;
    _T_1709_im <= _T_1708_im;
    _T_1710_re <= _T_1709_re;
    _T_1710_im <= _T_1709_im;
    _T_1711_re <= _T_1710_re;
    _T_1711_im <= _T_1710_im;
    _T_1712_re <= _T_1711_re;
    _T_1712_im <= _T_1711_im;
    _T_1713_re <= _T_1712_re;
    _T_1713_im <= _T_1712_im;
    _T_1714_re <= _T_1713_re;
    _T_1714_im <= _T_1713_im;
    _T_1715_re <= _T_1714_re;
    _T_1715_im <= _T_1714_im;
    _T_1716_re <= _T_1715_re;
    _T_1716_im <= _T_1715_im;
    _T_1717_re <= _T_1716_re;
    _T_1717_im <= _T_1716_im;
    _T_1718_re <= _T_1717_re;
    _T_1718_im <= _T_1717_im;
    _T_1719_re <= _T_1718_re;
    _T_1719_im <= _T_1718_im;
    _T_1720_re <= _T_1719_re;
    _T_1720_im <= _T_1719_im;
    _T_1721_re <= _T_1720_re;
    _T_1721_im <= _T_1720_im;
    _T_1722_re <= _T_1721_re;
    _T_1722_im <= _T_1721_im;
    _T_1723_re <= _T_1722_re;
    _T_1723_im <= _T_1722_im;
    _T_1724_re <= _T_1723_re;
    _T_1724_im <= _T_1723_im;
    _T_1725_re <= _T_1724_re;
    _T_1725_im <= _T_1724_im;
    _T_1726_re <= _T_1725_re;
    _T_1726_im <= _T_1725_im;
    _T_1727_re <= _T_1726_re;
    _T_1727_im <= _T_1726_im;
    _T_1728_re <= _T_1727_re;
    _T_1728_im <= _T_1727_im;
    _T_1729_re <= _T_1728_re;
    _T_1729_im <= _T_1728_im;
    _T_1730_re <= _T_1729_re;
    _T_1730_im <= _T_1729_im;
    _T_1731_re <= _T_1730_re;
    _T_1731_im <= _T_1730_im;
    _T_1732_re <= _T_1731_re;
    _T_1732_im <= _T_1731_im;
    _T_1733_re <= _T_1732_re;
    _T_1733_im <= _T_1732_im;
    _T_1734_re <= _T_1733_re;
    _T_1734_im <= _T_1733_im;
    _T_1735_re <= _T_1734_re;
    _T_1735_im <= _T_1734_im;
    _T_1736_re <= _T_1735_re;
    _T_1736_im <= _T_1735_im;
    _T_1737_re <= _T_1736_re;
    _T_1737_im <= _T_1736_im;
    _T_1738_re <= _T_1737_re;
    _T_1738_im <= _T_1737_im;
    _T_1739_re <= _T_1738_re;
    _T_1739_im <= _T_1738_im;
    _T_1740_re <= _T_1739_re;
    _T_1740_im <= _T_1739_im;
    _T_1741_re <= _T_1740_re;
    _T_1741_im <= _T_1740_im;
    _T_1742_re <= _T_1741_re;
    _T_1742_im <= _T_1741_im;
    _T_1743_re <= _T_1742_re;
    _T_1743_im <= _T_1742_im;
    _T_1744_re <= _T_1743_re;
    _T_1744_im <= _T_1743_im;
    _T_1745_re <= _T_1744_re;
    _T_1745_im <= _T_1744_im;
    _T_1746_re <= _T_1745_re;
    _T_1746_im <= _T_1745_im;
    _T_1747_re <= _T_1746_re;
    _T_1747_im <= _T_1746_im;
    _T_1748_re <= _T_1747_re;
    _T_1748_im <= _T_1747_im;
    _T_1749_re <= _T_1748_re;
    _T_1749_im <= _T_1748_im;
    _T_1750_re <= _T_1749_re;
    _T_1750_im <= _T_1749_im;
    _T_1751_re <= _T_1750_re;
    _T_1751_im <= _T_1750_im;
    _T_1752_re <= _T_1751_re;
    _T_1752_im <= _T_1751_im;
    _T_1753_re <= _T_1752_re;
    _T_1753_im <= _T_1752_im;
    _T_1754_re <= _T_1753_re;
    _T_1754_im <= _T_1753_im;
    _T_1755_re <= _T_1754_re;
    _T_1755_im <= _T_1754_im;
    _T_1756_re <= _T_1755_re;
    _T_1756_im <= _T_1755_im;
    _T_1757_re <= _T_1756_re;
    _T_1757_im <= _T_1756_im;
    _T_1758_re <= _T_1757_re;
    _T_1758_im <= _T_1757_im;
    _T_1759_re <= _T_1758_re;
    _T_1759_im <= _T_1758_im;
    _T_1760_re <= _T_1759_re;
    _T_1760_im <= _T_1759_im;
    _T_1761_re <= _T_1760_re;
    _T_1761_im <= _T_1760_im;
    _T_1762_re <= _T_1761_re;
    _T_1762_im <= _T_1761_im;
    _T_1763_re <= _T_1762_re;
    _T_1763_im <= _T_1762_im;
    _T_1764_re <= _T_1763_re;
    _T_1764_im <= _T_1763_im;
    _T_1765_re <= _T_1764_re;
    _T_1765_im <= _T_1764_im;
    _T_1766_re <= _T_1765_re;
    _T_1766_im <= _T_1765_im;
    _T_1767_re <= _T_1766_re;
    _T_1767_im <= _T_1766_im;
    _T_1768_re <= _T_1767_re;
    _T_1768_im <= _T_1767_im;
    _T_1769_re <= _T_1768_re;
    _T_1769_im <= _T_1768_im;
    _T_1770_re <= _T_1769_re;
    _T_1770_im <= _T_1769_im;
    _T_1771_re <= _T_1770_re;
    _T_1771_im <= _T_1770_im;
    _T_1772_re <= _T_1771_re;
    _T_1772_im <= _T_1771_im;
    _T_1773_re <= _T_1772_re;
    _T_1773_im <= _T_1772_im;
    _T_1774_re <= _T_1773_re;
    _T_1774_im <= _T_1773_im;
    _T_1775_re <= _T_1774_re;
    _T_1775_im <= _T_1774_im;
    _T_1776_re <= _T_1775_re;
    _T_1776_im <= _T_1775_im;
    _T_1777_re <= _T_1776_re;
    _T_1777_im <= _T_1776_im;
    _T_1778_re <= _T_1777_re;
    _T_1778_im <= _T_1777_im;
    _T_1779_re <= _T_1778_re;
    _T_1779_im <= _T_1778_im;
    _T_1780_re <= _T_1779_re;
    _T_1780_im <= _T_1779_im;
    _T_1781_re <= _T_1780_re;
    _T_1781_im <= _T_1780_im;
    _T_1782_re <= _T_1781_re;
    _T_1782_im <= _T_1781_im;
    _T_1783_re <= _T_1782_re;
    _T_1783_im <= _T_1782_im;
    _T_1784_re <= _T_1783_re;
    _T_1784_im <= _T_1783_im;
    _T_1785_re <= _T_1784_re;
    _T_1785_im <= _T_1784_im;
    _T_1786_re <= _T_1785_re;
    _T_1786_im <= _T_1785_im;
    _T_1787_re <= _T_1786_re;
    _T_1787_im <= _T_1786_im;
    _T_1788_re <= _T_1787_re;
    _T_1788_im <= _T_1787_im;
    _T_1789_re <= _T_1788_re;
    _T_1789_im <= _T_1788_im;
    _T_1790_re <= _T_1789_re;
    _T_1790_im <= _T_1789_im;
    _T_1791_re <= _T_1790_re;
    _T_1791_im <= _T_1790_im;
    _T_1792_re <= _T_1791_re;
    _T_1792_im <= _T_1791_im;
    _T_1793_re <= _T_1792_re;
    _T_1793_im <= _T_1792_im;
    _T_1794_re <= _T_1793_re;
    _T_1794_im <= _T_1793_im;
    _T_1795_re <= _T_1794_re;
    _T_1795_im <= _T_1794_im;
    _T_1796_re <= _T_1795_re;
    _T_1796_im <= _T_1795_im;
    _T_1797_re <= _T_1796_re;
    _T_1797_im <= _T_1796_im;
    _T_1798_re <= _T_1797_re;
    _T_1798_im <= _T_1797_im;
    _T_1799_re <= _T_1798_re;
    _T_1799_im <= _T_1798_im;
    _T_1800_re <= _T_1799_re;
    _T_1800_im <= _T_1799_im;
    _T_1801_re <= _T_1800_re;
    _T_1801_im <= _T_1800_im;
    _T_1802_re <= _T_1801_re;
    _T_1802_im <= _T_1801_im;
    _T_1803_re <= _T_1802_re;
    _T_1803_im <= _T_1802_im;
    _T_1804_re <= _T_1803_re;
    _T_1804_im <= _T_1803_im;
    _T_1805_re <= _T_1804_re;
    _T_1805_im <= _T_1804_im;
    _T_1806_re <= _T_1805_re;
    _T_1806_im <= _T_1805_im;
    _T_1807_re <= _T_1806_re;
    _T_1807_im <= _T_1806_im;
    _T_1808_re <= _T_1807_re;
    _T_1808_im <= _T_1807_im;
    _T_1809_re <= _T_1808_re;
    _T_1809_im <= _T_1808_im;
    _T_1810_re <= _T_1809_re;
    _T_1810_im <= _T_1809_im;
    _T_1811_re <= _T_1810_re;
    _T_1811_im <= _T_1810_im;
    _T_1812_re <= _T_1811_re;
    _T_1812_im <= _T_1811_im;
    _T_1813_re <= _T_1812_re;
    _T_1813_im <= _T_1812_im;
    _T_1814_re <= _T_1813_re;
    _T_1814_im <= _T_1813_im;
    _T_1815_re <= _T_1814_re;
    _T_1815_im <= _T_1814_im;
    _T_1816_re <= _T_1815_re;
    _T_1816_im <= _T_1815_im;
    _T_1817_re <= _T_1816_re;
    _T_1817_im <= _T_1816_im;
    _T_1818_re <= _T_1817_re;
    _T_1818_im <= _T_1817_im;
    _T_1819_re <= _T_1818_re;
    _T_1819_im <= _T_1818_im;
    _T_1820_re <= _T_1819_re;
    _T_1820_im <= _T_1819_im;
    _T_1821_re <= _T_1820_re;
    _T_1821_im <= _T_1820_im;
    _T_1822_re <= _T_1821_re;
    _T_1822_im <= _T_1821_im;
    _T_1823_re <= _T_1822_re;
    _T_1823_im <= _T_1822_im;
    _T_1824_re <= _T_1823_re;
    _T_1824_im <= _T_1823_im;
    _T_1825_re <= _T_1824_re;
    _T_1825_im <= _T_1824_im;
    _T_1826_re <= _T_1825_re;
    _T_1826_im <= _T_1825_im;
    _T_1827_re <= _T_1826_re;
    _T_1827_im <= _T_1826_im;
    _T_1828_re <= _T_1827_re;
    _T_1828_im <= _T_1827_im;
    _T_1829_re <= _T_1828_re;
    _T_1829_im <= _T_1828_im;
    _T_1830_re <= _T_1829_re;
    _T_1830_im <= _T_1829_im;
    _T_1831_re <= _T_1830_re;
    _T_1831_im <= _T_1830_im;
    _T_1832_re <= _T_1831_re;
    _T_1832_im <= _T_1831_im;
    _T_1833_re <= _T_1832_re;
    _T_1833_im <= _T_1832_im;
    _T_1834_re <= _T_1833_re;
    _T_1834_im <= _T_1833_im;
    _T_1835_re <= _T_1834_re;
    _T_1835_im <= _T_1834_im;
    _T_1836_re <= _T_1835_re;
    _T_1836_im <= _T_1835_im;
    _T_1837_re <= _T_1836_re;
    _T_1837_im <= _T_1836_im;
    _T_1838_re <= _T_1837_re;
    _T_1838_im <= _T_1837_im;
    _T_1839_re <= _T_1838_re;
    _T_1839_im <= _T_1838_im;
    _T_1840_re <= _T_1839_re;
    _T_1840_im <= _T_1839_im;
    _T_1841_re <= _T_1840_re;
    _T_1841_im <= _T_1840_im;
    _T_1842_re <= _T_1841_re;
    _T_1842_im <= _T_1841_im;
    _T_1843_re <= _T_1842_re;
    _T_1843_im <= _T_1842_im;
    _T_1844_re <= _T_1843_re;
    _T_1844_im <= _T_1843_im;
    _T_1845_re <= _T_1844_re;
    _T_1845_im <= _T_1844_im;
    _T_1846_re <= _T_1845_re;
    _T_1846_im <= _T_1845_im;
    _T_1847_re <= _T_1846_re;
    _T_1847_im <= _T_1846_im;
    _T_1848_re <= _T_1847_re;
    _T_1848_im <= _T_1847_im;
    _T_1849_re <= _T_1848_re;
    _T_1849_im <= _T_1848_im;
    _T_1850_re <= _T_1849_re;
    _T_1850_im <= _T_1849_im;
    _T_1851_re <= _T_1850_re;
    _T_1851_im <= _T_1850_im;
    _T_1852_re <= _T_1851_re;
    _T_1852_im <= _T_1851_im;
    _T_1853_re <= _T_1852_re;
    _T_1853_im <= _T_1852_im;
    _T_1854_re <= _T_1853_re;
    _T_1854_im <= _T_1853_im;
    _T_1855_re <= _T_1854_re;
    _T_1855_im <= _T_1854_im;
    _T_1856_re <= _T_1855_re;
    _T_1856_im <= _T_1855_im;
    _T_1857_re <= _T_1856_re;
    _T_1857_im <= _T_1856_im;
    _T_1858_re <= _T_1857_re;
    _T_1858_im <= _T_1857_im;
    _T_1859_re <= _T_1858_re;
    _T_1859_im <= _T_1858_im;
    _T_1860_re <= _T_1859_re;
    _T_1860_im <= _T_1859_im;
    _T_1861_re <= _T_1860_re;
    _T_1861_im <= _T_1860_im;
    _T_1862_re <= _T_1861_re;
    _T_1862_im <= _T_1861_im;
    _T_1863_re <= _T_1862_re;
    _T_1863_im <= _T_1862_im;
    _T_1864_re <= _T_1863_re;
    _T_1864_im <= _T_1863_im;
    _T_1865_re <= _T_1864_re;
    _T_1865_im <= _T_1864_im;
    _T_1866_re <= _T_1865_re;
    _T_1866_im <= _T_1865_im;
    _T_1867_re <= _T_1866_re;
    _T_1867_im <= _T_1866_im;
    _T_1868_re <= _T_1867_re;
    _T_1868_im <= _T_1867_im;
    _T_1869_re <= _T_1868_re;
    _T_1869_im <= _T_1868_im;
    _T_1870_re <= _T_1869_re;
    _T_1870_im <= _T_1869_im;
    _T_1871_re <= _T_1870_re;
    _T_1871_im <= _T_1870_im;
    _T_1872_re <= _T_1871_re;
    _T_1872_im <= _T_1871_im;
    _T_1873_re <= _T_1872_re;
    _T_1873_im <= _T_1872_im;
    _T_1874_re <= _T_1873_re;
    _T_1874_im <= _T_1873_im;
    _T_1875_re <= _T_1874_re;
    _T_1875_im <= _T_1874_im;
    _T_1876_re <= _T_1875_re;
    _T_1876_im <= _T_1875_im;
    _T_1877_re <= _T_1876_re;
    _T_1877_im <= _T_1876_im;
    _T_1878_re <= _T_1877_re;
    _T_1878_im <= _T_1877_im;
    _T_1879_re <= _T_1878_re;
    _T_1879_im <= _T_1878_im;
    _T_1880_re <= _T_1879_re;
    _T_1880_im <= _T_1879_im;
    _T_1881_re <= _T_1880_re;
    _T_1881_im <= _T_1880_im;
    _T_1882_re <= _T_1881_re;
    _T_1882_im <= _T_1881_im;
    _T_1883_re <= _T_1882_re;
    _T_1883_im <= _T_1882_im;
    _T_1884_re <= _T_1883_re;
    _T_1884_im <= _T_1883_im;
    _T_1885_re <= _T_1884_re;
    _T_1885_im <= _T_1884_im;
    _T_1886_re <= _T_1885_re;
    _T_1886_im <= _T_1885_im;
    _T_1887_re <= _T_1886_re;
    _T_1887_im <= _T_1886_im;
    _T_1888_re <= _T_1887_re;
    _T_1888_im <= _T_1887_im;
    _T_1889_re <= _T_1888_re;
    _T_1889_im <= _T_1888_im;
    _T_1890_re <= _T_1889_re;
    _T_1890_im <= _T_1889_im;
    _T_1891_re <= _T_1890_re;
    _T_1891_im <= _T_1890_im;
    _T_1892_re <= _T_1891_re;
    _T_1892_im <= _T_1891_im;
    _T_1893_re <= _T_1892_re;
    _T_1893_im <= _T_1892_im;
    _T_1894_re <= _T_1893_re;
    _T_1894_im <= _T_1893_im;
    _T_1895_re <= _T_1894_re;
    _T_1895_im <= _T_1894_im;
    _T_1896_re <= _T_1895_re;
    _T_1896_im <= _T_1895_im;
    _T_1897_re <= _T_1896_re;
    _T_1897_im <= _T_1896_im;
    _T_1898_re <= _T_1897_re;
    _T_1898_im <= _T_1897_im;
    _T_1899_re <= _T_1898_re;
    _T_1899_im <= _T_1898_im;
    _T_1900_re <= _T_1899_re;
    _T_1900_im <= _T_1899_im;
    _T_1901_re <= _T_1900_re;
    _T_1901_im <= _T_1900_im;
    _T_1902_re <= _T_1901_re;
    _T_1902_im <= _T_1901_im;
    _T_1903_re <= _T_1902_re;
    _T_1903_im <= _T_1902_im;
    _T_1904_re <= _T_1903_re;
    _T_1904_im <= _T_1903_im;
    _T_1905_re <= _T_1904_re;
    _T_1905_im <= _T_1904_im;
    _T_1906_re <= _T_1905_re;
    _T_1906_im <= _T_1905_im;
    _T_1907_re <= _T_1906_re;
    _T_1907_im <= _T_1906_im;
    _T_1908_re <= _T_1907_re;
    _T_1908_im <= _T_1907_im;
    _T_1909_re <= _T_1908_re;
    _T_1909_im <= _T_1908_im;
    _T_1910_re <= _T_1909_re;
    _T_1910_im <= _T_1909_im;
    _T_1911_re <= _T_1910_re;
    _T_1911_im <= _T_1910_im;
    _T_1912_re <= _T_1911_re;
    _T_1912_im <= _T_1911_im;
    _T_1913_re <= _T_1912_re;
    _T_1913_im <= _T_1912_im;
    _T_1914_re <= _T_1913_re;
    _T_1914_im <= _T_1913_im;
    _T_1915_re <= _T_1914_re;
    _T_1915_im <= _T_1914_im;
    _T_1916_re <= _T_1915_re;
    _T_1916_im <= _T_1915_im;
    _T_1917_re <= _T_1916_re;
    _T_1917_im <= _T_1916_im;
    _T_1918_re <= _T_1917_re;
    _T_1918_im <= _T_1917_im;
    _T_1919_re <= _T_1918_re;
    _T_1919_im <= _T_1918_im;
    _T_1920_re <= _T_1919_re;
    _T_1920_im <= _T_1919_im;
    _T_1921_re <= _T_1920_re;
    _T_1921_im <= _T_1920_im;
    _T_1922_re <= _T_1921_re;
    _T_1922_im <= _T_1921_im;
    _T_1923_re <= _T_1922_re;
    _T_1923_im <= _T_1922_im;
    _T_1924_re <= _T_1923_re;
    _T_1924_im <= _T_1923_im;
    _T_1925_re <= _T_1924_re;
    _T_1925_im <= _T_1924_im;
    _T_1926_re <= _T_1925_re;
    _T_1926_im <= _T_1925_im;
    _T_1927_re <= _T_1926_re;
    _T_1927_im <= _T_1926_im;
    _T_1928_re <= _T_1927_re;
    _T_1928_im <= _T_1927_im;
    _T_1929_re <= _T_1928_re;
    _T_1929_im <= _T_1928_im;
    _T_1930_re <= _T_1929_re;
    _T_1930_im <= _T_1929_im;
    _T_1931_re <= _T_1930_re;
    _T_1931_im <= _T_1930_im;
    _T_1932_re <= _T_1931_re;
    _T_1932_im <= _T_1931_im;
    _T_1933_re <= _T_1932_re;
    _T_1933_im <= _T_1932_im;
    _T_1934_re <= _T_1933_re;
    _T_1934_im <= _T_1933_im;
    _T_1935_re <= _T_1934_re;
    _T_1935_im <= _T_1934_im;
    _T_1936_re <= _T_1935_re;
    _T_1936_im <= _T_1935_im;
    _T_1937_re <= _T_1936_re;
    _T_1937_im <= _T_1936_im;
    _T_1938_re <= _T_1937_re;
    _T_1938_im <= _T_1937_im;
    _T_1939_re <= _T_1938_re;
    _T_1939_im <= _T_1938_im;
    _T_1940_re <= _T_1939_re;
    _T_1940_im <= _T_1939_im;
    _T_1941_re <= _T_1940_re;
    _T_1941_im <= _T_1940_im;
    _T_1942_re <= _T_1941_re;
    _T_1942_im <= _T_1941_im;
    _T_1943_re <= _T_1942_re;
    _T_1943_im <= _T_1942_im;
    _T_1944_re <= _T_1943_re;
    _T_1944_im <= _T_1943_im;
    _T_1945_re <= _T_1944_re;
    _T_1945_im <= _T_1944_im;
    _T_1946_re <= _T_1945_re;
    _T_1946_im <= _T_1945_im;
    _T_1947_re <= _T_1946_re;
    _T_1947_im <= _T_1946_im;
    _T_1948_re <= _T_1947_re;
    _T_1948_im <= _T_1947_im;
    _T_1949_re <= _T_1948_re;
    _T_1949_im <= _T_1948_im;
    _T_1950_re <= _T_1949_re;
    _T_1950_im <= _T_1949_im;
    _T_1951_re <= _T_1950_re;
    _T_1951_im <= _T_1950_im;
    _T_1952_re <= _T_1951_re;
    _T_1952_im <= _T_1951_im;
    _T_1953_re <= _T_1952_re;
    _T_1953_im <= _T_1952_im;
    _T_1954_re <= _T_1953_re;
    _T_1954_im <= _T_1953_im;
    _T_1955_re <= _T_1954_re;
    _T_1955_im <= _T_1954_im;
    _T_1956_re <= _T_1955_re;
    _T_1956_im <= _T_1955_im;
    _T_1957_re <= _T_1956_re;
    _T_1957_im <= _T_1956_im;
    _T_1958_re <= _T_1957_re;
    _T_1958_im <= _T_1957_im;
    _T_1959_re <= _T_1958_re;
    _T_1959_im <= _T_1958_im;
    _T_1960_re <= _T_1959_re;
    _T_1960_im <= _T_1959_im;
    _T_1961_re <= _T_1960_re;
    _T_1961_im <= _T_1960_im;
    _T_1962_re <= _T_1961_re;
    _T_1962_im <= _T_1961_im;
    _T_1963_re <= _T_1962_re;
    _T_1963_im <= _T_1962_im;
    _T_1964_re <= _T_1963_re;
    _T_1964_im <= _T_1963_im;
    _T_1965_re <= _T_1964_re;
    _T_1965_im <= _T_1964_im;
    _T_1966_re <= _T_1965_re;
    _T_1966_im <= _T_1965_im;
    _T_1967_re <= _T_1966_re;
    _T_1967_im <= _T_1966_im;
    _T_1968_re <= _T_1967_re;
    _T_1968_im <= _T_1967_im;
    _T_1969_re <= _T_1968_re;
    _T_1969_im <= _T_1968_im;
    _T_1970_re <= _T_1969_re;
    _T_1970_im <= _T_1969_im;
    _T_1971_re <= _T_1970_re;
    _T_1971_im <= _T_1970_im;
    _T_1972_re <= _T_1971_re;
    _T_1972_im <= _T_1971_im;
    _T_1973_re <= _T_1972_re;
    _T_1973_im <= _T_1972_im;
    _T_1974_re <= _T_1973_re;
    _T_1974_im <= _T_1973_im;
    _T_1975_re <= _T_1974_re;
    _T_1975_im <= _T_1974_im;
    _T_1976_re <= _T_1975_re;
    _T_1976_im <= _T_1975_im;
    _T_1977_re <= _T_1976_re;
    _T_1977_im <= _T_1976_im;
    _T_1978_re <= _T_1977_re;
    _T_1978_im <= _T_1977_im;
    _T_1979_re <= _T_1978_re;
    _T_1979_im <= _T_1978_im;
    _T_1980_re <= _T_1979_re;
    _T_1980_im <= _T_1979_im;
    _T_1981_re <= _T_1980_re;
    _T_1981_im <= _T_1980_im;
    _T_1982_re <= _T_1981_re;
    _T_1982_im <= _T_1981_im;
    _T_1983_re <= _T_1982_re;
    _T_1983_im <= _T_1982_im;
    _T_1984_re <= _T_1983_re;
    _T_1984_im <= _T_1983_im;
    _T_1985_re <= _T_1984_re;
    _T_1985_im <= _T_1984_im;
    _T_1986_re <= _T_1985_re;
    _T_1986_im <= _T_1985_im;
    _T_1987_re <= _T_1986_re;
    _T_1987_im <= _T_1986_im;
    _T_1988_re <= _T_1987_re;
    _T_1988_im <= _T_1987_im;
    _T_1989_re <= _T_1988_re;
    _T_1989_im <= _T_1988_im;
    _T_1990_re <= _T_1989_re;
    _T_1990_im <= _T_1989_im;
    _T_1991_re <= _T_1990_re;
    _T_1991_im <= _T_1990_im;
    _T_1992_re <= _T_1991_re;
    _T_1992_im <= _T_1991_im;
    _T_1993_re <= _T_1992_re;
    _T_1993_im <= _T_1992_im;
    _T_1994_re <= _T_1993_re;
    _T_1994_im <= _T_1993_im;
    _T_1995_re <= _T_1994_re;
    _T_1995_im <= _T_1994_im;
    _T_1996_re <= _T_1995_re;
    _T_1996_im <= _T_1995_im;
    _T_1997_re <= _T_1996_re;
    _T_1997_im <= _T_1996_im;
    _T_1998_re <= _T_1997_re;
    _T_1998_im <= _T_1997_im;
    _T_1999_re <= _T_1998_re;
    _T_1999_im <= _T_1998_im;
    _T_2000_re <= _T_1999_re;
    _T_2000_im <= _T_1999_im;
    _T_2001_re <= _T_2000_re;
    _T_2001_im <= _T_2000_im;
    _T_2002_re <= _T_2001_re;
    _T_2002_im <= _T_2001_im;
    _T_2003_re <= _T_2002_re;
    _T_2003_im <= _T_2002_im;
    _T_2004_re <= _T_2003_re;
    _T_2004_im <= _T_2003_im;
    _T_2005_re <= _T_2004_re;
    _T_2005_im <= _T_2004_im;
    _T_2006_re <= _T_2005_re;
    _T_2006_im <= _T_2005_im;
    _T_2007_re <= _T_2006_re;
    _T_2007_im <= _T_2006_im;
    _T_2008_re <= _T_2007_re;
    _T_2008_im <= _T_2007_im;
    _T_2009_re <= _T_2008_re;
    _T_2009_im <= _T_2008_im;
    _T_2010_re <= _T_2009_re;
    _T_2010_im <= _T_2009_im;
    _T_2011_re <= _T_2010_re;
    _T_2011_im <= _T_2010_im;
    _T_2012_re <= _T_2011_re;
    _T_2012_im <= _T_2011_im;
    _T_2013_re <= _T_2012_re;
    _T_2013_im <= _T_2012_im;
    _T_2014_re <= _T_2013_re;
    _T_2014_im <= _T_2013_im;
    _T_2015_re <= _T_2014_re;
    _T_2015_im <= _T_2014_im;
    _T_2016_re <= _T_2015_re;
    _T_2016_im <= _T_2015_im;
    _T_2017_re <= _T_2016_re;
    _T_2017_im <= _T_2016_im;
    _T_2018_re <= _T_2017_re;
    _T_2018_im <= _T_2017_im;
    _T_2019_re <= _T_2018_re;
    _T_2019_im <= _T_2018_im;
    _T_2020_re <= _T_2019_re;
    _T_2020_im <= _T_2019_im;
    _T_2021_re <= _T_2020_re;
    _T_2021_im <= _T_2020_im;
    _T_2022_re <= _T_2021_re;
    _T_2022_im <= _T_2021_im;
    _T_2023_re <= _T_2022_re;
    _T_2023_im <= _T_2022_im;
    _T_2024_re <= _T_2023_re;
    _T_2024_im <= _T_2023_im;
    _T_2025_re <= _T_2024_re;
    _T_2025_im <= _T_2024_im;
    _T_2026_re <= _T_2025_re;
    _T_2026_im <= _T_2025_im;
    _T_2027_re <= _T_2026_re;
    _T_2027_im <= _T_2026_im;
    _T_2028_re <= _T_2027_re;
    _T_2028_im <= _T_2027_im;
    _T_2029_re <= _T_2028_re;
    _T_2029_im <= _T_2028_im;
    _T_2030_re <= _T_2029_re;
    _T_2030_im <= _T_2029_im;
    _T_2031_re <= _T_2030_re;
    _T_2031_im <= _T_2030_im;
    _T_2032_re <= _T_2031_re;
    _T_2032_im <= _T_2031_im;
    _T_2033_re <= _T_2032_re;
    _T_2033_im <= _T_2032_im;
    _T_2034_re <= _T_2033_re;
    _T_2034_im <= _T_2033_im;
    _T_2035_re <= _T_2034_re;
    _T_2035_im <= _T_2034_im;
    _T_2036_re <= _T_2035_re;
    _T_2036_im <= _T_2035_im;
    _T_2037_re <= _T_2036_re;
    _T_2037_im <= _T_2036_im;
    _T_2038_re <= _T_2037_re;
    _T_2038_im <= _T_2037_im;
    _T_2039_re <= _T_2038_re;
    _T_2039_im <= _T_2038_im;
    _T_2040_re <= _T_2039_re;
    _T_2040_im <= _T_2039_im;
    _T_2041_re <= _T_2040_re;
    _T_2041_im <= _T_2040_im;
    _T_2042_re <= _T_2041_re;
    _T_2042_im <= _T_2041_im;
    _T_2043_re <= _T_2042_re;
    _T_2043_im <= _T_2042_im;
    _T_2044_re <= _T_2043_re;
    _T_2044_im <= _T_2043_im;
    _T_2045_re <= _T_2044_re;
    _T_2045_im <= _T_2044_im;
    _T_2046_re <= _T_2045_re;
    _T_2046_im <= _T_2045_im;
    _T_2047_re <= _T_2046_re;
    _T_2047_im <= _T_2046_im;
    _T_2048_re <= _T_2047_re;
    _T_2048_im <= _T_2047_im;
    _T_2049_re <= _T_2048_re;
    _T_2049_im <= _T_2048_im;
    _T_2050_re <= _T_2049_re;
    _T_2050_im <= _T_2049_im;
    _T_2051_re <= _T_2050_re;
    _T_2051_im <= _T_2050_im;
    _T_2052_re <= _T_2051_re;
    _T_2052_im <= _T_2051_im;
    _T_2053_re <= _T_2052_re;
    _T_2053_im <= _T_2052_im;
    _T_2054_re <= _T_2053_re;
    _T_2054_im <= _T_2053_im;
    _T_2055_re <= _T_2054_re;
    _T_2055_im <= _T_2054_im;
    _T_2056_re <= _T_2055_re;
    _T_2056_im <= _T_2055_im;
    _T_2057_re <= _T_2056_re;
    _T_2057_im <= _T_2056_im;
    _T_2058_re <= _T_2057_re;
    _T_2058_im <= _T_2057_im;
    _T_2059_re <= _T_2058_re;
    _T_2059_im <= _T_2058_im;
    _T_2060_re <= _T_2059_re;
    _T_2060_im <= _T_2059_im;
    _T_2061_re <= _T_2060_re;
    _T_2061_im <= _T_2060_im;
    _T_2062_re <= _T_2061_re;
    _T_2062_im <= _T_2061_im;
    _T_2063_re <= _T_2062_re;
    _T_2063_im <= _T_2062_im;
    _T_2064_re <= _T_2063_re;
    _T_2064_im <= _T_2063_im;
    _T_2065_re <= _T_2064_re;
    _T_2065_im <= _T_2064_im;
    _T_2066_re <= _T_2065_re;
    _T_2066_im <= _T_2065_im;
    _T_2067_re <= _T_2066_re;
    _T_2067_im <= _T_2066_im;
    _T_2068_re <= _T_2067_re;
    _T_2068_im <= _T_2067_im;
    _T_2069_re <= _T_2068_re;
    _T_2069_im <= _T_2068_im;
    _T_2070_re <= _T_2069_re;
    _T_2070_im <= _T_2069_im;
    _T_2071_re <= _T_2070_re;
    _T_2071_im <= _T_2070_im;
    _T_2072_re <= _T_2071_re;
    _T_2072_im <= _T_2071_im;
    _T_2073_re <= _T_2072_re;
    _T_2073_im <= _T_2072_im;
    _T_2074_re <= _T_2073_re;
    _T_2074_im <= _T_2073_im;
    _T_2075_re <= _T_2074_re;
    _T_2075_im <= _T_2074_im;
    _T_2076_re <= _T_2075_re;
    _T_2076_im <= _T_2075_im;
    _T_2077_re <= _T_2076_re;
    _T_2077_im <= _T_2076_im;
    _T_2078_re <= _T_2077_re;
    _T_2078_im <= _T_2077_im;
    _T_2079_re <= _T_2078_re;
    _T_2079_im <= _T_2078_im;
    _T_2080_re <= _T_2079_re;
    _T_2080_im <= _T_2079_im;
    _T_2081_re <= _T_2080_re;
    _T_2081_im <= _T_2080_im;
    _T_2082_re <= _T_2081_re;
    _T_2082_im <= _T_2081_im;
    _T_2083_re <= _T_2082_re;
    _T_2083_im <= _T_2082_im;
    _T_2084_re <= _T_2083_re;
    _T_2084_im <= _T_2083_im;
    _T_2085_re <= _T_2084_re;
    _T_2085_im <= _T_2084_im;
    _T_2086_re <= _T_2085_re;
    _T_2086_im <= _T_2085_im;
    _T_2087_re <= _T_2086_re;
    _T_2087_im <= _T_2086_im;
    _T_2088_re <= _T_2087_re;
    _T_2088_im <= _T_2087_im;
    _T_2089_re <= _T_2088_re;
    _T_2089_im <= _T_2088_im;
    _T_2090_re <= _T_2089_re;
    _T_2090_im <= _T_2089_im;
    _T_2091_re <= _T_2090_re;
    _T_2091_im <= _T_2090_im;
    _T_2092_re <= _T_2091_re;
    _T_2092_im <= _T_2091_im;
    _T_2093_re <= _T_2092_re;
    _T_2093_im <= _T_2092_im;
    _T_2094_re <= _T_2093_re;
    _T_2094_im <= _T_2093_im;
    _T_2095_re <= _T_2094_re;
    _T_2095_im <= _T_2094_im;
    _T_2096_re <= _T_2095_re;
    _T_2096_im <= _T_2095_im;
    _T_2097_re <= _T_2096_re;
    _T_2097_im <= _T_2096_im;
    _T_2098_re <= _T_2097_re;
    _T_2098_im <= _T_2097_im;
    _T_2099_re <= _T_2098_re;
    _T_2099_im <= _T_2098_im;
    _T_2100_re <= _T_2099_re;
    _T_2100_im <= _T_2099_im;
    _T_2101_re <= _T_2100_re;
    _T_2101_im <= _T_2100_im;
    _T_2102_re <= _T_2101_re;
    _T_2102_im <= _T_2101_im;
    _T_2103_re <= _T_2102_re;
    _T_2103_im <= _T_2102_im;
    _T_2104_re <= _T_2103_re;
    _T_2104_im <= _T_2103_im;
    _T_2105_re <= _T_2104_re;
    _T_2105_im <= _T_2104_im;
    _T_2106_re <= _T_2105_re;
    _T_2106_im <= _T_2105_im;
    _T_2107_re <= _T_2106_re;
    _T_2107_im <= _T_2106_im;
    _T_2108_re <= _T_2107_re;
    _T_2108_im <= _T_2107_im;
    _T_2109_re <= _T_2108_re;
    _T_2109_im <= _T_2108_im;
    _T_2110_re <= _T_2109_re;
    _T_2110_im <= _T_2109_im;
    _T_2111_re <= _T_2110_re;
    _T_2111_im <= _T_2110_im;
    _T_2112_re <= _T_2111_re;
    _T_2112_im <= _T_2111_im;
    _T_2113_re <= _T_2112_re;
    _T_2113_im <= _T_2112_im;
    _T_2114_re <= _T_2113_re;
    _T_2114_im <= _T_2113_im;
    _T_2115_re <= _T_2114_re;
    _T_2115_im <= _T_2114_im;
    _T_2116_re <= _T_2115_re;
    _T_2116_im <= _T_2115_im;
    _T_2117_re <= _T_2116_re;
    _T_2117_im <= _T_2116_im;
    _T_2118_re <= _T_2117_re;
    _T_2118_im <= _T_2117_im;
    _T_2119_re <= _T_2118_re;
    _T_2119_im <= _T_2118_im;
    _T_2120_re <= _T_2119_re;
    _T_2120_im <= _T_2119_im;
    _T_2121_re <= _T_2120_re;
    _T_2121_im <= _T_2120_im;
    _T_2122_re <= _T_2121_re;
    _T_2122_im <= _T_2121_im;
    _T_2123_re <= _T_2122_re;
    _T_2123_im <= _T_2122_im;
    _T_2124_re <= _T_2123_re;
    _T_2124_im <= _T_2123_im;
    _T_2125_re <= _T_2124_re;
    _T_2125_im <= _T_2124_im;
    _T_2126_re <= _T_2125_re;
    _T_2126_im <= _T_2125_im;
    _T_2127_re <= _T_2126_re;
    _T_2127_im <= _T_2126_im;
    _T_2128_re <= _T_2127_re;
    _T_2128_im <= _T_2127_im;
    _T_2129_re <= _T_2128_re;
    _T_2129_im <= _T_2128_im;
    _T_2130_re <= _T_2129_re;
    _T_2130_im <= _T_2129_im;
    _T_2131_re <= _T_2130_re;
    _T_2131_im <= _T_2130_im;
    _T_2132_re <= _T_2131_re;
    _T_2132_im <= _T_2131_im;
    _T_2133_re <= _T_2132_re;
    _T_2133_im <= _T_2132_im;
    _T_2134_re <= _T_2133_re;
    _T_2134_im <= _T_2133_im;
    _T_2135_re <= _T_2134_re;
    _T_2135_im <= _T_2134_im;
    _T_2136_re <= _T_2135_re;
    _T_2136_im <= _T_2135_im;
    _T_2137_re <= _T_2136_re;
    _T_2137_im <= _T_2136_im;
    _T_2138_re <= _T_2137_re;
    _T_2138_im <= _T_2137_im;
    _T_2139_re <= _T_2138_re;
    _T_2139_im <= _T_2138_im;
    _T_2140_re <= _T_2139_re;
    _T_2140_im <= _T_2139_im;
    _T_2141_re <= _T_2140_re;
    _T_2141_im <= _T_2140_im;
    _T_2142_re <= _T_2141_re;
    _T_2142_im <= _T_2141_im;
    _T_2143_re <= _T_2142_re;
    _T_2143_im <= _T_2142_im;
    _T_2144_re <= _T_2143_re;
    _T_2144_im <= _T_2143_im;
    _T_2145_re <= _T_2144_re;
    _T_2145_im <= _T_2144_im;
    _T_2146_re <= _T_2145_re;
    _T_2146_im <= _T_2145_im;
    _T_2147_re <= _T_2146_re;
    _T_2147_im <= _T_2146_im;
    _T_2148_re <= _T_2147_re;
    _T_2148_im <= _T_2147_im;
    _T_2149_re <= _T_2148_re;
    _T_2149_im <= _T_2148_im;
    _T_2150_re <= _T_2149_re;
    _T_2150_im <= _T_2149_im;
    _T_2151_re <= _T_2150_re;
    _T_2151_im <= _T_2150_im;
    _T_2152_re <= _T_2151_re;
    _T_2152_im <= _T_2151_im;
    _T_2153_re <= _T_2152_re;
    _T_2153_im <= _T_2152_im;
    _T_2154_re <= _T_2153_re;
    _T_2154_im <= _T_2153_im;
    _T_2155_re <= _T_2154_re;
    _T_2155_im <= _T_2154_im;
    _T_2156_re <= _T_2155_re;
    _T_2156_im <= _T_2155_im;
    _T_2157_re <= _T_2156_re;
    _T_2157_im <= _T_2156_im;
    _T_2158_re <= _T_2157_re;
    _T_2158_im <= _T_2157_im;
    _T_2159_re <= _T_2158_re;
    _T_2159_im <= _T_2158_im;
    _T_2160_re <= _T_2159_re;
    _T_2160_im <= _T_2159_im;
    _T_2161_re <= _T_2160_re;
    _T_2161_im <= _T_2160_im;
    _T_2162_re <= _T_2161_re;
    _T_2162_im <= _T_2161_im;
    _T_2163_re <= _T_2162_re;
    _T_2163_im <= _T_2162_im;
    _T_2164_re <= _T_2163_re;
    _T_2164_im <= _T_2163_im;
    _T_2165_re <= _T_2164_re;
    _T_2165_im <= _T_2164_im;
    _T_2166_re <= _T_2165_re;
    _T_2166_im <= _T_2165_im;
    _T_2167_re <= _T_2166_re;
    _T_2167_im <= _T_2166_im;
    _T_2168_re <= _T_2167_re;
    _T_2168_im <= _T_2167_im;
    _T_2169_re <= _T_2168_re;
    _T_2169_im <= _T_2168_im;
    _T_2170_re <= _T_2169_re;
    _T_2170_im <= _T_2169_im;
    _T_2171_re <= _T_2170_re;
    _T_2171_im <= _T_2170_im;
    _T_2172_re <= _T_2171_re;
    _T_2172_im <= _T_2171_im;
    _T_2173_re <= _T_2172_re;
    _T_2173_im <= _T_2172_im;
    _T_2174_re <= _T_2173_re;
    _T_2174_im <= _T_2173_im;
    _T_2175_re <= _T_2174_re;
    _T_2175_im <= _T_2174_im;
    _T_2176_re <= _T_2175_re;
    _T_2176_im <= _T_2175_im;
    _T_2177_re <= _T_2176_re;
    _T_2177_im <= _T_2176_im;
    _T_2178_re <= _T_2177_re;
    _T_2178_im <= _T_2177_im;
    _T_2179_re <= _T_2178_re;
    _T_2179_im <= _T_2178_im;
    _T_2180_re <= _T_2179_re;
    _T_2180_im <= _T_2179_im;
    _T_2181_re <= _T_2180_re;
    _T_2181_im <= _T_2180_im;
    _T_2182_re <= _T_2181_re;
    _T_2182_im <= _T_2181_im;
    _T_2183_re <= _T_2182_re;
    _T_2183_im <= _T_2182_im;
    _T_2184_re <= _T_2183_re;
    _T_2184_im <= _T_2183_im;
    _T_2185_re <= _T_2184_re;
    _T_2185_im <= _T_2184_im;
    _T_2186_re <= _T_2185_re;
    _T_2186_im <= _T_2185_im;
    _T_2187_re <= _T_2186_re;
    _T_2187_im <= _T_2186_im;
    _T_2188_re <= _T_2187_re;
    _T_2188_im <= _T_2187_im;
    _T_2189_re <= _T_2188_re;
    _T_2189_im <= _T_2188_im;
    _T_2190_re <= _T_2189_re;
    _T_2190_im <= _T_2189_im;
    _T_2191_re <= _T_2190_re;
    _T_2191_im <= _T_2190_im;
    _T_2192_re <= _T_2191_re;
    _T_2192_im <= _T_2191_im;
    _T_2193_re <= _T_2192_re;
    _T_2193_im <= _T_2192_im;
    _T_2194_re <= _T_2193_re;
    _T_2194_im <= _T_2193_im;
    _T_2195_re <= _T_2194_re;
    _T_2195_im <= _T_2194_im;
    _T_2196_re <= _T_2195_re;
    _T_2196_im <= _T_2195_im;
    _T_2197_re <= _T_2196_re;
    _T_2197_im <= _T_2196_im;
    _T_2198_re <= _T_2197_re;
    _T_2198_im <= _T_2197_im;
    _T_2199_re <= _T_2198_re;
    _T_2199_im <= _T_2198_im;
    _T_2200_re <= _T_2199_re;
    _T_2200_im <= _T_2199_im;
    _T_2201_re <= _T_2200_re;
    _T_2201_im <= _T_2200_im;
    _T_2202_re <= _T_2201_re;
    _T_2202_im <= _T_2201_im;
    _T_2203_re <= _T_2202_re;
    _T_2203_im <= _T_2202_im;
    _T_2204_re <= _T_2203_re;
    _T_2204_im <= _T_2203_im;
    _T_2205_re <= _T_2204_re;
    _T_2205_im <= _T_2204_im;
    _T_2206_re <= _T_2205_re;
    _T_2206_im <= _T_2205_im;
    _T_2207_re <= _T_2206_re;
    _T_2207_im <= _T_2206_im;
    _T_2208_re <= _T_2207_re;
    _T_2208_im <= _T_2207_im;
    _T_2209_re <= _T_2208_re;
    _T_2209_im <= _T_2208_im;
    _T_2210_re <= _T_2209_re;
    _T_2210_im <= _T_2209_im;
    _T_2211_re <= _T_2210_re;
    _T_2211_im <= _T_2210_im;
    _T_2212_re <= _T_2211_re;
    _T_2212_im <= _T_2211_im;
    _T_2213_re <= _T_2212_re;
    _T_2213_im <= _T_2212_im;
    _T_2214_re <= _T_2213_re;
    _T_2214_im <= _T_2213_im;
    _T_2215_re <= _T_2214_re;
    _T_2215_im <= _T_2214_im;
    _T_2216_re <= _T_2215_re;
    _T_2216_im <= _T_2215_im;
    _T_2217_re <= _T_2216_re;
    _T_2217_im <= _T_2216_im;
    _T_2218_re <= _T_2217_re;
    _T_2218_im <= _T_2217_im;
    _T_2219_re <= _T_2218_re;
    _T_2219_im <= _T_2218_im;
    _T_2220_re <= _T_2219_re;
    _T_2220_im <= _T_2219_im;
    _T_2221_re <= _T_2220_re;
    _T_2221_im <= _T_2220_im;
    _T_2222_re <= _T_2221_re;
    _T_2222_im <= _T_2221_im;
    _T_2223_re <= _T_2222_re;
    _T_2223_im <= _T_2222_im;
    _T_2224_re <= _T_2223_re;
    _T_2224_im <= _T_2223_im;
    _T_2225_re <= _T_2224_re;
    _T_2225_im <= _T_2224_im;
    _T_2226_re <= _T_2225_re;
    _T_2226_im <= _T_2225_im;
    _T_2227_re <= _T_2226_re;
    _T_2227_im <= _T_2226_im;
    _T_2228_re <= _T_2227_re;
    _T_2228_im <= _T_2227_im;
    _T_2229_re <= _T_2228_re;
    _T_2229_im <= _T_2228_im;
    _T_2230_re <= _T_2229_re;
    _T_2230_im <= _T_2229_im;
    _T_2231_re <= _T_2230_re;
    _T_2231_im <= _T_2230_im;
    _T_2232_re <= _T_2231_re;
    _T_2232_im <= _T_2231_im;
    _T_2233_re <= _T_2232_re;
    _T_2233_im <= _T_2232_im;
    _T_2234_re <= _T_2233_re;
    _T_2234_im <= _T_2233_im;
    _T_2235_re <= _T_2234_re;
    _T_2235_im <= _T_2234_im;
    _T_2236_re <= _T_2235_re;
    _T_2236_im <= _T_2235_im;
    _T_2239_re <= Butterfly_io_out2_re;
    _T_2239_im <= Butterfly_io_out2_im;
    _T_2240_re <= _T_2239_re;
    _T_2240_im <= _T_2239_im;
    _T_2241_re <= _T_2240_re;
    _T_2241_im <= _T_2240_im;
    _T_2242_re <= _T_2241_re;
    _T_2242_im <= _T_2241_im;
    _T_2243_re <= _T_2242_re;
    _T_2243_im <= _T_2242_im;
    _T_2244_re <= _T_2243_re;
    _T_2244_im <= _T_2243_im;
    _T_2245_re <= _T_2244_re;
    _T_2245_im <= _T_2244_im;
    _T_2246_re <= _T_2245_re;
    _T_2246_im <= _T_2245_im;
    _T_2247_re <= _T_2246_re;
    _T_2247_im <= _T_2246_im;
    _T_2248_re <= _T_2247_re;
    _T_2248_im <= _T_2247_im;
    _T_2249_re <= _T_2248_re;
    _T_2249_im <= _T_2248_im;
    _T_2250_re <= _T_2249_re;
    _T_2250_im <= _T_2249_im;
    _T_2251_re <= _T_2250_re;
    _T_2251_im <= _T_2250_im;
    _T_2252_re <= _T_2251_re;
    _T_2252_im <= _T_2251_im;
    _T_2253_re <= _T_2252_re;
    _T_2253_im <= _T_2252_im;
    _T_2254_re <= _T_2253_re;
    _T_2254_im <= _T_2253_im;
    _T_2255_re <= _T_2254_re;
    _T_2255_im <= _T_2254_im;
    _T_2256_re <= _T_2255_re;
    _T_2256_im <= _T_2255_im;
    _T_2257_re <= _T_2256_re;
    _T_2257_im <= _T_2256_im;
    _T_2258_re <= _T_2257_re;
    _T_2258_im <= _T_2257_im;
    _T_2259_re <= _T_2258_re;
    _T_2259_im <= _T_2258_im;
    _T_2260_re <= _T_2259_re;
    _T_2260_im <= _T_2259_im;
    _T_2261_re <= _T_2260_re;
    _T_2261_im <= _T_2260_im;
    _T_2262_re <= _T_2261_re;
    _T_2262_im <= _T_2261_im;
    _T_2263_re <= _T_2262_re;
    _T_2263_im <= _T_2262_im;
    _T_2264_re <= _T_2263_re;
    _T_2264_im <= _T_2263_im;
    _T_2265_re <= _T_2264_re;
    _T_2265_im <= _T_2264_im;
    _T_2266_re <= _T_2265_re;
    _T_2266_im <= _T_2265_im;
    _T_2267_re <= _T_2266_re;
    _T_2267_im <= _T_2266_im;
    _T_2268_re <= _T_2267_re;
    _T_2268_im <= _T_2267_im;
    _T_2269_re <= _T_2268_re;
    _T_2269_im <= _T_2268_im;
    _T_2270_re <= _T_2269_re;
    _T_2270_im <= _T_2269_im;
    _T_2271_re <= _T_2270_re;
    _T_2271_im <= _T_2270_im;
    _T_2272_re <= _T_2271_re;
    _T_2272_im <= _T_2271_im;
    _T_2273_re <= _T_2272_re;
    _T_2273_im <= _T_2272_im;
    _T_2274_re <= _T_2273_re;
    _T_2274_im <= _T_2273_im;
    _T_2275_re <= _T_2274_re;
    _T_2275_im <= _T_2274_im;
    _T_2276_re <= _T_2275_re;
    _T_2276_im <= _T_2275_im;
    _T_2277_re <= _T_2276_re;
    _T_2277_im <= _T_2276_im;
    _T_2278_re <= _T_2277_re;
    _T_2278_im <= _T_2277_im;
    _T_2279_re <= _T_2278_re;
    _T_2279_im <= _T_2278_im;
    _T_2280_re <= _T_2279_re;
    _T_2280_im <= _T_2279_im;
    _T_2281_re <= _T_2280_re;
    _T_2281_im <= _T_2280_im;
    _T_2282_re <= _T_2281_re;
    _T_2282_im <= _T_2281_im;
    _T_2283_re <= _T_2282_re;
    _T_2283_im <= _T_2282_im;
    _T_2284_re <= _T_2283_re;
    _T_2284_im <= _T_2283_im;
    _T_2285_re <= _T_2284_re;
    _T_2285_im <= _T_2284_im;
    _T_2286_re <= _T_2285_re;
    _T_2286_im <= _T_2285_im;
    _T_2287_re <= _T_2286_re;
    _T_2287_im <= _T_2286_im;
    _T_2288_re <= _T_2287_re;
    _T_2288_im <= _T_2287_im;
    _T_2289_re <= _T_2288_re;
    _T_2289_im <= _T_2288_im;
    _T_2290_re <= _T_2289_re;
    _T_2290_im <= _T_2289_im;
    _T_2291_re <= _T_2290_re;
    _T_2291_im <= _T_2290_im;
    _T_2292_re <= _T_2291_re;
    _T_2292_im <= _T_2291_im;
    _T_2293_re <= _T_2292_re;
    _T_2293_im <= _T_2292_im;
    _T_2294_re <= _T_2293_re;
    _T_2294_im <= _T_2293_im;
    _T_2295_re <= _T_2294_re;
    _T_2295_im <= _T_2294_im;
    _T_2296_re <= _T_2295_re;
    _T_2296_im <= _T_2295_im;
    _T_2297_re <= _T_2296_re;
    _T_2297_im <= _T_2296_im;
    _T_2298_re <= _T_2297_re;
    _T_2298_im <= _T_2297_im;
    _T_2299_re <= _T_2298_re;
    _T_2299_im <= _T_2298_im;
    _T_2300_re <= _T_2299_re;
    _T_2300_im <= _T_2299_im;
    _T_2301_re <= _T_2300_re;
    _T_2301_im <= _T_2300_im;
    _T_2302_re <= _T_2301_re;
    _T_2302_im <= _T_2301_im;
    _T_2303_re <= _T_2302_re;
    _T_2303_im <= _T_2302_im;
    _T_2304_re <= _T_2303_re;
    _T_2304_im <= _T_2303_im;
    _T_2305_re <= _T_2304_re;
    _T_2305_im <= _T_2304_im;
    _T_2306_re <= _T_2305_re;
    _T_2306_im <= _T_2305_im;
    _T_2307_re <= _T_2306_re;
    _T_2307_im <= _T_2306_im;
    _T_2308_re <= _T_2307_re;
    _T_2308_im <= _T_2307_im;
    _T_2309_re <= _T_2308_re;
    _T_2309_im <= _T_2308_im;
    _T_2310_re <= _T_2309_re;
    _T_2310_im <= _T_2309_im;
    _T_2311_re <= _T_2310_re;
    _T_2311_im <= _T_2310_im;
    _T_2312_re <= _T_2311_re;
    _T_2312_im <= _T_2311_im;
    _T_2313_re <= _T_2312_re;
    _T_2313_im <= _T_2312_im;
    _T_2314_re <= _T_2313_re;
    _T_2314_im <= _T_2313_im;
    _T_2315_re <= _T_2314_re;
    _T_2315_im <= _T_2314_im;
    _T_2316_re <= _T_2315_re;
    _T_2316_im <= _T_2315_im;
    _T_2317_re <= _T_2316_re;
    _T_2317_im <= _T_2316_im;
    _T_2318_re <= _T_2317_re;
    _T_2318_im <= _T_2317_im;
    _T_2319_re <= _T_2318_re;
    _T_2319_im <= _T_2318_im;
    _T_2320_re <= _T_2319_re;
    _T_2320_im <= _T_2319_im;
    _T_2321_re <= _T_2320_re;
    _T_2321_im <= _T_2320_im;
    _T_2322_re <= _T_2321_re;
    _T_2322_im <= _T_2321_im;
    _T_2323_re <= _T_2322_re;
    _T_2323_im <= _T_2322_im;
    _T_2324_re <= _T_2323_re;
    _T_2324_im <= _T_2323_im;
    _T_2325_re <= _T_2324_re;
    _T_2325_im <= _T_2324_im;
    _T_2326_re <= _T_2325_re;
    _T_2326_im <= _T_2325_im;
    _T_2327_re <= _T_2326_re;
    _T_2327_im <= _T_2326_im;
    _T_2328_re <= _T_2327_re;
    _T_2328_im <= _T_2327_im;
    _T_2329_re <= _T_2328_re;
    _T_2329_im <= _T_2328_im;
    _T_2330_re <= _T_2329_re;
    _T_2330_im <= _T_2329_im;
    _T_2331_re <= _T_2330_re;
    _T_2331_im <= _T_2330_im;
    _T_2332_re <= _T_2331_re;
    _T_2332_im <= _T_2331_im;
    _T_2333_re <= _T_2332_re;
    _T_2333_im <= _T_2332_im;
    _T_2334_re <= _T_2333_re;
    _T_2334_im <= _T_2333_im;
    _T_2335_re <= _T_2334_re;
    _T_2335_im <= _T_2334_im;
    _T_2336_re <= _T_2335_re;
    _T_2336_im <= _T_2335_im;
    _T_2337_re <= _T_2336_re;
    _T_2337_im <= _T_2336_im;
    _T_2338_re <= _T_2337_re;
    _T_2338_im <= _T_2337_im;
    _T_2339_re <= _T_2338_re;
    _T_2339_im <= _T_2338_im;
    _T_2340_re <= _T_2339_re;
    _T_2340_im <= _T_2339_im;
    _T_2341_re <= _T_2340_re;
    _T_2341_im <= _T_2340_im;
    _T_2342_re <= _T_2341_re;
    _T_2342_im <= _T_2341_im;
    _T_2343_re <= _T_2342_re;
    _T_2343_im <= _T_2342_im;
    _T_2344_re <= _T_2343_re;
    _T_2344_im <= _T_2343_im;
    _T_2345_re <= _T_2344_re;
    _T_2345_im <= _T_2344_im;
    _T_2346_re <= _T_2345_re;
    _T_2346_im <= _T_2345_im;
    _T_2347_re <= _T_2346_re;
    _T_2347_im <= _T_2346_im;
    _T_2348_re <= _T_2347_re;
    _T_2348_im <= _T_2347_im;
    _T_2349_re <= _T_2348_re;
    _T_2349_im <= _T_2348_im;
    _T_2350_re <= _T_2349_re;
    _T_2350_im <= _T_2349_im;
    _T_2351_re <= _T_2350_re;
    _T_2351_im <= _T_2350_im;
    _T_2352_re <= _T_2351_re;
    _T_2352_im <= _T_2351_im;
    _T_2353_re <= _T_2352_re;
    _T_2353_im <= _T_2352_im;
    _T_2354_re <= _T_2353_re;
    _T_2354_im <= _T_2353_im;
    _T_2355_re <= _T_2354_re;
    _T_2355_im <= _T_2354_im;
    _T_2356_re <= _T_2355_re;
    _T_2356_im <= _T_2355_im;
    _T_2357_re <= _T_2356_re;
    _T_2357_im <= _T_2356_im;
    _T_2358_re <= _T_2357_re;
    _T_2358_im <= _T_2357_im;
    _T_2359_re <= _T_2358_re;
    _T_2359_im <= _T_2358_im;
    _T_2360_re <= _T_2359_re;
    _T_2360_im <= _T_2359_im;
    _T_2361_re <= _T_2360_re;
    _T_2361_im <= _T_2360_im;
    _T_2362_re <= _T_2361_re;
    _T_2362_im <= _T_2361_im;
    _T_2363_re <= _T_2362_re;
    _T_2363_im <= _T_2362_im;
    _T_2364_re <= _T_2363_re;
    _T_2364_im <= _T_2363_im;
    _T_2365_re <= _T_2364_re;
    _T_2365_im <= _T_2364_im;
    _T_2366_re <= _T_2365_re;
    _T_2366_im <= _T_2365_im;
    _T_2367_re <= _T_2366_re;
    _T_2367_im <= _T_2366_im;
    _T_2368_re <= _T_2367_re;
    _T_2368_im <= _T_2367_im;
    _T_2369_re <= _T_2368_re;
    _T_2369_im <= _T_2368_im;
    _T_2370_re <= _T_2369_re;
    _T_2370_im <= _T_2369_im;
    _T_2371_re <= _T_2370_re;
    _T_2371_im <= _T_2370_im;
    _T_2372_re <= _T_2371_re;
    _T_2372_im <= _T_2371_im;
    _T_2373_re <= _T_2372_re;
    _T_2373_im <= _T_2372_im;
    _T_2374_re <= _T_2373_re;
    _T_2374_im <= _T_2373_im;
    _T_2375_re <= _T_2374_re;
    _T_2375_im <= _T_2374_im;
    _T_2376_re <= _T_2375_re;
    _T_2376_im <= _T_2375_im;
    _T_2377_re <= _T_2376_re;
    _T_2377_im <= _T_2376_im;
    _T_2378_re <= _T_2377_re;
    _T_2378_im <= _T_2377_im;
    _T_2379_re <= _T_2378_re;
    _T_2379_im <= _T_2378_im;
    _T_2380_re <= _T_2379_re;
    _T_2380_im <= _T_2379_im;
    _T_2381_re <= _T_2380_re;
    _T_2381_im <= _T_2380_im;
    _T_2382_re <= _T_2381_re;
    _T_2382_im <= _T_2381_im;
    _T_2383_re <= _T_2382_re;
    _T_2383_im <= _T_2382_im;
    _T_2384_re <= _T_2383_re;
    _T_2384_im <= _T_2383_im;
    _T_2385_re <= _T_2384_re;
    _T_2385_im <= _T_2384_im;
    _T_2386_re <= _T_2385_re;
    _T_2386_im <= _T_2385_im;
    _T_2387_re <= _T_2386_re;
    _T_2387_im <= _T_2386_im;
    _T_2388_re <= _T_2387_re;
    _T_2388_im <= _T_2387_im;
    _T_2389_re <= _T_2388_re;
    _T_2389_im <= _T_2388_im;
    _T_2390_re <= _T_2389_re;
    _T_2390_im <= _T_2389_im;
    _T_2391_re <= _T_2390_re;
    _T_2391_im <= _T_2390_im;
    _T_2392_re <= _T_2391_re;
    _T_2392_im <= _T_2391_im;
    _T_2393_re <= _T_2392_re;
    _T_2393_im <= _T_2392_im;
    _T_2394_re <= _T_2393_re;
    _T_2394_im <= _T_2393_im;
    _T_2395_re <= _T_2394_re;
    _T_2395_im <= _T_2394_im;
    _T_2396_re <= _T_2395_re;
    _T_2396_im <= _T_2395_im;
    _T_2397_re <= _T_2396_re;
    _T_2397_im <= _T_2396_im;
    _T_2398_re <= _T_2397_re;
    _T_2398_im <= _T_2397_im;
    _T_2399_re <= _T_2398_re;
    _T_2399_im <= _T_2398_im;
    _T_2400_re <= _T_2399_re;
    _T_2400_im <= _T_2399_im;
    _T_2401_re <= _T_2400_re;
    _T_2401_im <= _T_2400_im;
    _T_2402_re <= _T_2401_re;
    _T_2402_im <= _T_2401_im;
    _T_2403_re <= _T_2402_re;
    _T_2403_im <= _T_2402_im;
    _T_2404_re <= _T_2403_re;
    _T_2404_im <= _T_2403_im;
    _T_2405_re <= _T_2404_re;
    _T_2405_im <= _T_2404_im;
    _T_2406_re <= _T_2405_re;
    _T_2406_im <= _T_2405_im;
    _T_2407_re <= _T_2406_re;
    _T_2407_im <= _T_2406_im;
    _T_2408_re <= _T_2407_re;
    _T_2408_im <= _T_2407_im;
    _T_2409_re <= _T_2408_re;
    _T_2409_im <= _T_2408_im;
    _T_2410_re <= _T_2409_re;
    _T_2410_im <= _T_2409_im;
    _T_2411_re <= _T_2410_re;
    _T_2411_im <= _T_2410_im;
    _T_2412_re <= _T_2411_re;
    _T_2412_im <= _T_2411_im;
    _T_2413_re <= _T_2412_re;
    _T_2413_im <= _T_2412_im;
    _T_2414_re <= _T_2413_re;
    _T_2414_im <= _T_2413_im;
    _T_2415_re <= _T_2414_re;
    _T_2415_im <= _T_2414_im;
    _T_2416_re <= _T_2415_re;
    _T_2416_im <= _T_2415_im;
    _T_2417_re <= _T_2416_re;
    _T_2417_im <= _T_2416_im;
    _T_2418_re <= _T_2417_re;
    _T_2418_im <= _T_2417_im;
    _T_2419_re <= _T_2418_re;
    _T_2419_im <= _T_2418_im;
    _T_2420_re <= _T_2419_re;
    _T_2420_im <= _T_2419_im;
    _T_2421_re <= _T_2420_re;
    _T_2421_im <= _T_2420_im;
    _T_2422_re <= _T_2421_re;
    _T_2422_im <= _T_2421_im;
    _T_2423_re <= _T_2422_re;
    _T_2423_im <= _T_2422_im;
    _T_2424_re <= _T_2423_re;
    _T_2424_im <= _T_2423_im;
    _T_2425_re <= _T_2424_re;
    _T_2425_im <= _T_2424_im;
    _T_2426_re <= _T_2425_re;
    _T_2426_im <= _T_2425_im;
    _T_2427_re <= _T_2426_re;
    _T_2427_im <= _T_2426_im;
    _T_2428_re <= _T_2427_re;
    _T_2428_im <= _T_2427_im;
    _T_2429_re <= _T_2428_re;
    _T_2429_im <= _T_2428_im;
    _T_2430_re <= _T_2429_re;
    _T_2430_im <= _T_2429_im;
    _T_2431_re <= _T_2430_re;
    _T_2431_im <= _T_2430_im;
    _T_2432_re <= _T_2431_re;
    _T_2432_im <= _T_2431_im;
    _T_2433_re <= _T_2432_re;
    _T_2433_im <= _T_2432_im;
    _T_2434_re <= _T_2433_re;
    _T_2434_im <= _T_2433_im;
    _T_2435_re <= _T_2434_re;
    _T_2435_im <= _T_2434_im;
    _T_2436_re <= _T_2435_re;
    _T_2436_im <= _T_2435_im;
    _T_2437_re <= _T_2436_re;
    _T_2437_im <= _T_2436_im;
    _T_2438_re <= _T_2437_re;
    _T_2438_im <= _T_2437_im;
    _T_2439_re <= _T_2438_re;
    _T_2439_im <= _T_2438_im;
    _T_2440_re <= _T_2439_re;
    _T_2440_im <= _T_2439_im;
    _T_2441_re <= _T_2440_re;
    _T_2441_im <= _T_2440_im;
    _T_2442_re <= _T_2441_re;
    _T_2442_im <= _T_2441_im;
    _T_2443_re <= _T_2442_re;
    _T_2443_im <= _T_2442_im;
    _T_2444_re <= _T_2443_re;
    _T_2444_im <= _T_2443_im;
    _T_2445_re <= _T_2444_re;
    _T_2445_im <= _T_2444_im;
    _T_2446_re <= _T_2445_re;
    _T_2446_im <= _T_2445_im;
    _T_2447_re <= _T_2446_re;
    _T_2447_im <= _T_2446_im;
    _T_2448_re <= _T_2447_re;
    _T_2448_im <= _T_2447_im;
    _T_2449_re <= _T_2448_re;
    _T_2449_im <= _T_2448_im;
    _T_2450_re <= _T_2449_re;
    _T_2450_im <= _T_2449_im;
    _T_2451_re <= _T_2450_re;
    _T_2451_im <= _T_2450_im;
    _T_2452_re <= _T_2451_re;
    _T_2452_im <= _T_2451_im;
    _T_2453_re <= _T_2452_re;
    _T_2453_im <= _T_2452_im;
    _T_2454_re <= _T_2453_re;
    _T_2454_im <= _T_2453_im;
    _T_2455_re <= _T_2454_re;
    _T_2455_im <= _T_2454_im;
    _T_2456_re <= _T_2455_re;
    _T_2456_im <= _T_2455_im;
    _T_2457_re <= _T_2456_re;
    _T_2457_im <= _T_2456_im;
    _T_2458_re <= _T_2457_re;
    _T_2458_im <= _T_2457_im;
    _T_2459_re <= _T_2458_re;
    _T_2459_im <= _T_2458_im;
    _T_2460_re <= _T_2459_re;
    _T_2460_im <= _T_2459_im;
    _T_2461_re <= _T_2460_re;
    _T_2461_im <= _T_2460_im;
    _T_2462_re <= _T_2461_re;
    _T_2462_im <= _T_2461_im;
    _T_2463_re <= _T_2462_re;
    _T_2463_im <= _T_2462_im;
    _T_2464_re <= _T_2463_re;
    _T_2464_im <= _T_2463_im;
    _T_2465_re <= _T_2464_re;
    _T_2465_im <= _T_2464_im;
    _T_2466_re <= _T_2465_re;
    _T_2466_im <= _T_2465_im;
    _T_2467_re <= _T_2466_re;
    _T_2467_im <= _T_2466_im;
    _T_2468_re <= _T_2467_re;
    _T_2468_im <= _T_2467_im;
    _T_2469_re <= _T_2468_re;
    _T_2469_im <= _T_2468_im;
    _T_2470_re <= _T_2469_re;
    _T_2470_im <= _T_2469_im;
    _T_2471_re <= _T_2470_re;
    _T_2471_im <= _T_2470_im;
    _T_2472_re <= _T_2471_re;
    _T_2472_im <= _T_2471_im;
    _T_2473_re <= _T_2472_re;
    _T_2473_im <= _T_2472_im;
    _T_2474_re <= _T_2473_re;
    _T_2474_im <= _T_2473_im;
    _T_2475_re <= _T_2474_re;
    _T_2475_im <= _T_2474_im;
    _T_2476_re <= _T_2475_re;
    _T_2476_im <= _T_2475_im;
    _T_2477_re <= _T_2476_re;
    _T_2477_im <= _T_2476_im;
    _T_2478_re <= _T_2477_re;
    _T_2478_im <= _T_2477_im;
    _T_2479_re <= _T_2478_re;
    _T_2479_im <= _T_2478_im;
    _T_2480_re <= _T_2479_re;
    _T_2480_im <= _T_2479_im;
    _T_2481_re <= _T_2480_re;
    _T_2481_im <= _T_2480_im;
    _T_2482_re <= _T_2481_re;
    _T_2482_im <= _T_2481_im;
    _T_2483_re <= _T_2482_re;
    _T_2483_im <= _T_2482_im;
    _T_2484_re <= _T_2483_re;
    _T_2484_im <= _T_2483_im;
    _T_2485_re <= _T_2484_re;
    _T_2485_im <= _T_2484_im;
    _T_2486_re <= _T_2485_re;
    _T_2486_im <= _T_2485_im;
    _T_2487_re <= _T_2486_re;
    _T_2487_im <= _T_2486_im;
    _T_2488_re <= _T_2487_re;
    _T_2488_im <= _T_2487_im;
    _T_2489_re <= _T_2488_re;
    _T_2489_im <= _T_2488_im;
    _T_2490_re <= _T_2489_re;
    _T_2490_im <= _T_2489_im;
    _T_2491_re <= _T_2490_re;
    _T_2491_im <= _T_2490_im;
    _T_2492_re <= _T_2491_re;
    _T_2492_im <= _T_2491_im;
    _T_2493_re <= _T_2492_re;
    _T_2493_im <= _T_2492_im;
    _T_2494_re <= _T_2493_re;
    _T_2494_im <= _T_2493_im;
    _T_2495_re <= _T_2494_re;
    _T_2495_im <= _T_2494_im;
    _T_2496_re <= _T_2495_re;
    _T_2496_im <= _T_2495_im;
    _T_2497_re <= _T_2496_re;
    _T_2497_im <= _T_2496_im;
    _T_2498_re <= _T_2497_re;
    _T_2498_im <= _T_2497_im;
    _T_2499_re <= _T_2498_re;
    _T_2499_im <= _T_2498_im;
    _T_2500_re <= _T_2499_re;
    _T_2500_im <= _T_2499_im;
    _T_2501_re <= _T_2500_re;
    _T_2501_im <= _T_2500_im;
    _T_2502_re <= _T_2501_re;
    _T_2502_im <= _T_2501_im;
    _T_2503_re <= _T_2502_re;
    _T_2503_im <= _T_2502_im;
    _T_2504_re <= _T_2503_re;
    _T_2504_im <= _T_2503_im;
    _T_2505_re <= _T_2504_re;
    _T_2505_im <= _T_2504_im;
    _T_2506_re <= _T_2505_re;
    _T_2506_im <= _T_2505_im;
    _T_2507_re <= _T_2506_re;
    _T_2507_im <= _T_2506_im;
    _T_2508_re <= _T_2507_re;
    _T_2508_im <= _T_2507_im;
    _T_2509_re <= _T_2508_re;
    _T_2509_im <= _T_2508_im;
    _T_2510_re <= _T_2509_re;
    _T_2510_im <= _T_2509_im;
    _T_2511_re <= _T_2510_re;
    _T_2511_im <= _T_2510_im;
    _T_2512_re <= _T_2511_re;
    _T_2512_im <= _T_2511_im;
    _T_2513_re <= _T_2512_re;
    _T_2513_im <= _T_2512_im;
    _T_2514_re <= _T_2513_re;
    _T_2514_im <= _T_2513_im;
    _T_2515_re <= _T_2514_re;
    _T_2515_im <= _T_2514_im;
    _T_2516_re <= _T_2515_re;
    _T_2516_im <= _T_2515_im;
    _T_2517_re <= _T_2516_re;
    _T_2517_im <= _T_2516_im;
    _T_2518_re <= _T_2517_re;
    _T_2518_im <= _T_2517_im;
    _T_2519_re <= _T_2518_re;
    _T_2519_im <= _T_2518_im;
    _T_2520_re <= _T_2519_re;
    _T_2520_im <= _T_2519_im;
    _T_2521_re <= _T_2520_re;
    _T_2521_im <= _T_2520_im;
    _T_2522_re <= _T_2521_re;
    _T_2522_im <= _T_2521_im;
    _T_2523_re <= _T_2522_re;
    _T_2523_im <= _T_2522_im;
    _T_2524_re <= _T_2523_re;
    _T_2524_im <= _T_2523_im;
    _T_2525_re <= _T_2524_re;
    _T_2525_im <= _T_2524_im;
    _T_2526_re <= _T_2525_re;
    _T_2526_im <= _T_2525_im;
    _T_2527_re <= _T_2526_re;
    _T_2527_im <= _T_2526_im;
    _T_2528_re <= _T_2527_re;
    _T_2528_im <= _T_2527_im;
    _T_2529_re <= _T_2528_re;
    _T_2529_im <= _T_2528_im;
    _T_2530_re <= _T_2529_re;
    _T_2530_im <= _T_2529_im;
    _T_2531_re <= _T_2530_re;
    _T_2531_im <= _T_2530_im;
    _T_2532_re <= _T_2531_re;
    _T_2532_im <= _T_2531_im;
    _T_2533_re <= _T_2532_re;
    _T_2533_im <= _T_2532_im;
    _T_2534_re <= _T_2533_re;
    _T_2534_im <= _T_2533_im;
    _T_2535_re <= _T_2534_re;
    _T_2535_im <= _T_2534_im;
    _T_2536_re <= _T_2535_re;
    _T_2536_im <= _T_2535_im;
    _T_2537_re <= _T_2536_re;
    _T_2537_im <= _T_2536_im;
    _T_2538_re <= _T_2537_re;
    _T_2538_im <= _T_2537_im;
    _T_2539_re <= _T_2538_re;
    _T_2539_im <= _T_2538_im;
    _T_2540_re <= _T_2539_re;
    _T_2540_im <= _T_2539_im;
    _T_2541_re <= _T_2540_re;
    _T_2541_im <= _T_2540_im;
    _T_2542_re <= _T_2541_re;
    _T_2542_im <= _T_2541_im;
    _T_2543_re <= _T_2542_re;
    _T_2543_im <= _T_2542_im;
    _T_2544_re <= _T_2543_re;
    _T_2544_im <= _T_2543_im;
    _T_2545_re <= _T_2544_re;
    _T_2545_im <= _T_2544_im;
    _T_2546_re <= _T_2545_re;
    _T_2546_im <= _T_2545_im;
    _T_2547_re <= _T_2546_re;
    _T_2547_im <= _T_2546_im;
    _T_2548_re <= _T_2547_re;
    _T_2548_im <= _T_2547_im;
    _T_2549_re <= _T_2548_re;
    _T_2549_im <= _T_2548_im;
    _T_2550_re <= _T_2549_re;
    _T_2550_im <= _T_2549_im;
    _T_2551_re <= _T_2550_re;
    _T_2551_im <= _T_2550_im;
    _T_2552_re <= _T_2551_re;
    _T_2552_im <= _T_2551_im;
    _T_2553_re <= _T_2552_re;
    _T_2553_im <= _T_2552_im;
    _T_2554_re <= _T_2553_re;
    _T_2554_im <= _T_2553_im;
    _T_2555_re <= _T_2554_re;
    _T_2555_im <= _T_2554_im;
    _T_2556_re <= _T_2555_re;
    _T_2556_im <= _T_2555_im;
    _T_2557_re <= _T_2556_re;
    _T_2557_im <= _T_2556_im;
    _T_2558_re <= _T_2557_re;
    _T_2558_im <= _T_2557_im;
    _T_2559_re <= _T_2558_re;
    _T_2559_im <= _T_2558_im;
    _T_2560_re <= _T_2559_re;
    _T_2560_im <= _T_2559_im;
    _T_2561_re <= _T_2560_re;
    _T_2561_im <= _T_2560_im;
    _T_2562_re <= _T_2561_re;
    _T_2562_im <= _T_2561_im;
    _T_2563_re <= _T_2562_re;
    _T_2563_im <= _T_2562_im;
    _T_2564_re <= _T_2563_re;
    _T_2564_im <= _T_2563_im;
    _T_2565_re <= _T_2564_re;
    _T_2565_im <= _T_2564_im;
    _T_2566_re <= _T_2565_re;
    _T_2566_im <= _T_2565_im;
    _T_2567_re <= _T_2566_re;
    _T_2567_im <= _T_2566_im;
    _T_2568_re <= _T_2567_re;
    _T_2568_im <= _T_2567_im;
    _T_2569_re <= _T_2568_re;
    _T_2569_im <= _T_2568_im;
    _T_2570_re <= _T_2569_re;
    _T_2570_im <= _T_2569_im;
    _T_2571_re <= _T_2570_re;
    _T_2571_im <= _T_2570_im;
    _T_2572_re <= _T_2571_re;
    _T_2572_im <= _T_2571_im;
    _T_2573_re <= _T_2572_re;
    _T_2573_im <= _T_2572_im;
    _T_2574_re <= _T_2573_re;
    _T_2574_im <= _T_2573_im;
    _T_2575_re <= _T_2574_re;
    _T_2575_im <= _T_2574_im;
    _T_2576_re <= _T_2575_re;
    _T_2576_im <= _T_2575_im;
    _T_2577_re <= _T_2576_re;
    _T_2577_im <= _T_2576_im;
    _T_2578_re <= _T_2577_re;
    _T_2578_im <= _T_2577_im;
    _T_2579_re <= _T_2578_re;
    _T_2579_im <= _T_2578_im;
    _T_2580_re <= _T_2579_re;
    _T_2580_im <= _T_2579_im;
    _T_2581_re <= _T_2580_re;
    _T_2581_im <= _T_2580_im;
    _T_2582_re <= _T_2581_re;
    _T_2582_im <= _T_2581_im;
    _T_2583_re <= _T_2582_re;
    _T_2583_im <= _T_2582_im;
    _T_2584_re <= _T_2583_re;
    _T_2584_im <= _T_2583_im;
    _T_2585_re <= _T_2584_re;
    _T_2585_im <= _T_2584_im;
    _T_2586_re <= _T_2585_re;
    _T_2586_im <= _T_2585_im;
    _T_2587_re <= _T_2586_re;
    _T_2587_im <= _T_2586_im;
    _T_2588_re <= _T_2587_re;
    _T_2588_im <= _T_2587_im;
    _T_2589_re <= _T_2588_re;
    _T_2589_im <= _T_2588_im;
    _T_2590_re <= _T_2589_re;
    _T_2590_im <= _T_2589_im;
    _T_2591_re <= _T_2590_re;
    _T_2591_im <= _T_2590_im;
    _T_2592_re <= _T_2591_re;
    _T_2592_im <= _T_2591_im;
    _T_2593_re <= _T_2592_re;
    _T_2593_im <= _T_2592_im;
    _T_2594_re <= _T_2593_re;
    _T_2594_im <= _T_2593_im;
    _T_2595_re <= _T_2594_re;
    _T_2595_im <= _T_2594_im;
    _T_2596_re <= _T_2595_re;
    _T_2596_im <= _T_2595_im;
    _T_2597_re <= _T_2596_re;
    _T_2597_im <= _T_2596_im;
    _T_2598_re <= _T_2597_re;
    _T_2598_im <= _T_2597_im;
    _T_2599_re <= _T_2598_re;
    _T_2599_im <= _T_2598_im;
    _T_2600_re <= _T_2599_re;
    _T_2600_im <= _T_2599_im;
    _T_2601_re <= _T_2600_re;
    _T_2601_im <= _T_2600_im;
    _T_2602_re <= _T_2601_re;
    _T_2602_im <= _T_2601_im;
    _T_2603_re <= _T_2602_re;
    _T_2603_im <= _T_2602_im;
    _T_2604_re <= _T_2603_re;
    _T_2604_im <= _T_2603_im;
    _T_2605_re <= _T_2604_re;
    _T_2605_im <= _T_2604_im;
    _T_2606_re <= _T_2605_re;
    _T_2606_im <= _T_2605_im;
    _T_2607_re <= _T_2606_re;
    _T_2607_im <= _T_2606_im;
    _T_2608_re <= _T_2607_re;
    _T_2608_im <= _T_2607_im;
    _T_2609_re <= _T_2608_re;
    _T_2609_im <= _T_2608_im;
    _T_2610_re <= _T_2609_re;
    _T_2610_im <= _T_2609_im;
    _T_2611_re <= _T_2610_re;
    _T_2611_im <= _T_2610_im;
    _T_2612_re <= _T_2611_re;
    _T_2612_im <= _T_2611_im;
    _T_2613_re <= _T_2612_re;
    _T_2613_im <= _T_2612_im;
    _T_2614_re <= _T_2613_re;
    _T_2614_im <= _T_2613_im;
    _T_2615_re <= _T_2614_re;
    _T_2615_im <= _T_2614_im;
    _T_2616_re <= _T_2615_re;
    _T_2616_im <= _T_2615_im;
    _T_2617_re <= _T_2616_re;
    _T_2617_im <= _T_2616_im;
    _T_2618_re <= _T_2617_re;
    _T_2618_im <= _T_2617_im;
    _T_2619_re <= _T_2618_re;
    _T_2619_im <= _T_2618_im;
    _T_2620_re <= _T_2619_re;
    _T_2620_im <= _T_2619_im;
    _T_2621_re <= _T_2620_re;
    _T_2621_im <= _T_2620_im;
    _T_2622_re <= _T_2621_re;
    _T_2622_im <= _T_2621_im;
    _T_2623_re <= _T_2622_re;
    _T_2623_im <= _T_2622_im;
    _T_2624_re <= _T_2623_re;
    _T_2624_im <= _T_2623_im;
    _T_2625_re <= _T_2624_re;
    _T_2625_im <= _T_2624_im;
    _T_2626_re <= _T_2625_re;
    _T_2626_im <= _T_2625_im;
    _T_2627_re <= _T_2626_re;
    _T_2627_im <= _T_2626_im;
    _T_2628_re <= _T_2627_re;
    _T_2628_im <= _T_2627_im;
    _T_2629_re <= _T_2628_re;
    _T_2629_im <= _T_2628_im;
    _T_2630_re <= _T_2629_re;
    _T_2630_im <= _T_2629_im;
    _T_2631_re <= _T_2630_re;
    _T_2631_im <= _T_2630_im;
    _T_2632_re <= _T_2631_re;
    _T_2632_im <= _T_2631_im;
    _T_2633_re <= _T_2632_re;
    _T_2633_im <= _T_2632_im;
    _T_2634_re <= _T_2633_re;
    _T_2634_im <= _T_2633_im;
    _T_2635_re <= _T_2634_re;
    _T_2635_im <= _T_2634_im;
    _T_2636_re <= _T_2635_re;
    _T_2636_im <= _T_2635_im;
    _T_2637_re <= _T_2636_re;
    _T_2637_im <= _T_2636_im;
    _T_2638_re <= _T_2637_re;
    _T_2638_im <= _T_2637_im;
    _T_2639_re <= _T_2638_re;
    _T_2639_im <= _T_2638_im;
    _T_2640_re <= _T_2639_re;
    _T_2640_im <= _T_2639_im;
    _T_2641_re <= _T_2640_re;
    _T_2641_im <= _T_2640_im;
    _T_2642_re <= _T_2641_re;
    _T_2642_im <= _T_2641_im;
    _T_2643_re <= _T_2642_re;
    _T_2643_im <= _T_2642_im;
    _T_2644_re <= _T_2643_re;
    _T_2644_im <= _T_2643_im;
    _T_2645_re <= _T_2644_re;
    _T_2645_im <= _T_2644_im;
    _T_2646_re <= _T_2645_re;
    _T_2646_im <= _T_2645_im;
    _T_2647_re <= _T_2646_re;
    _T_2647_im <= _T_2646_im;
    _T_2648_re <= _T_2647_re;
    _T_2648_im <= _T_2647_im;
    _T_2649_re <= _T_2648_re;
    _T_2649_im <= _T_2648_im;
    _T_2650_re <= _T_2649_re;
    _T_2650_im <= _T_2649_im;
    _T_2651_re <= _T_2650_re;
    _T_2651_im <= _T_2650_im;
    _T_2652_re <= _T_2651_re;
    _T_2652_im <= _T_2651_im;
    _T_2653_re <= _T_2652_re;
    _T_2653_im <= _T_2652_im;
    _T_2654_re <= _T_2653_re;
    _T_2654_im <= _T_2653_im;
    _T_2655_re <= _T_2654_re;
    _T_2655_im <= _T_2654_im;
    _T_2656_re <= _T_2655_re;
    _T_2656_im <= _T_2655_im;
    _T_2657_re <= _T_2656_re;
    _T_2657_im <= _T_2656_im;
    _T_2658_re <= _T_2657_re;
    _T_2658_im <= _T_2657_im;
    _T_2659_re <= _T_2658_re;
    _T_2659_im <= _T_2658_im;
    _T_2660_re <= _T_2659_re;
    _T_2660_im <= _T_2659_im;
    _T_2661_re <= _T_2660_re;
    _T_2661_im <= _T_2660_im;
    _T_2662_re <= _T_2661_re;
    _T_2662_im <= _T_2661_im;
    _T_2663_re <= _T_2662_re;
    _T_2663_im <= _T_2662_im;
    _T_2664_re <= _T_2663_re;
    _T_2664_im <= _T_2663_im;
    _T_2665_re <= _T_2664_re;
    _T_2665_im <= _T_2664_im;
    _T_2666_re <= _T_2665_re;
    _T_2666_im <= _T_2665_im;
    _T_2667_re <= _T_2666_re;
    _T_2667_im <= _T_2666_im;
    _T_2668_re <= _T_2667_re;
    _T_2668_im <= _T_2667_im;
    _T_2669_re <= _T_2668_re;
    _T_2669_im <= _T_2668_im;
    _T_2670_re <= _T_2669_re;
    _T_2670_im <= _T_2669_im;
    _T_2671_re <= _T_2670_re;
    _T_2671_im <= _T_2670_im;
    _T_2672_re <= _T_2671_re;
    _T_2672_im <= _T_2671_im;
    _T_2673_re <= _T_2672_re;
    _T_2673_im <= _T_2672_im;
    _T_2674_re <= _T_2673_re;
    _T_2674_im <= _T_2673_im;
    _T_2675_re <= _T_2674_re;
    _T_2675_im <= _T_2674_im;
    _T_2676_re <= _T_2675_re;
    _T_2676_im <= _T_2675_im;
    _T_2677_re <= _T_2676_re;
    _T_2677_im <= _T_2676_im;
    _T_2678_re <= _T_2677_re;
    _T_2678_im <= _T_2677_im;
    _T_2679_re <= _T_2678_re;
    _T_2679_im <= _T_2678_im;
    _T_2680_re <= _T_2679_re;
    _T_2680_im <= _T_2679_im;
    _T_2681_re <= _T_2680_re;
    _T_2681_im <= _T_2680_im;
    _T_2682_re <= _T_2681_re;
    _T_2682_im <= _T_2681_im;
    _T_2683_re <= _T_2682_re;
    _T_2683_im <= _T_2682_im;
    _T_2684_re <= _T_2683_re;
    _T_2684_im <= _T_2683_im;
    _T_2685_re <= _T_2684_re;
    _T_2685_im <= _T_2684_im;
    _T_2686_re <= _T_2685_re;
    _T_2686_im <= _T_2685_im;
    _T_2687_re <= _T_2686_re;
    _T_2687_im <= _T_2686_im;
    _T_2688_re <= _T_2687_re;
    _T_2688_im <= _T_2687_im;
    _T_2689_re <= _T_2688_re;
    _T_2689_im <= _T_2688_im;
    _T_2690_re <= _T_2689_re;
    _T_2690_im <= _T_2689_im;
    _T_2691_re <= _T_2690_re;
    _T_2691_im <= _T_2690_im;
    _T_2692_re <= _T_2691_re;
    _T_2692_im <= _T_2691_im;
    _T_2693_re <= _T_2692_re;
    _T_2693_im <= _T_2692_im;
    _T_2694_re <= _T_2693_re;
    _T_2694_im <= _T_2693_im;
    _T_2695_re <= _T_2694_re;
    _T_2695_im <= _T_2694_im;
    _T_2696_re <= _T_2695_re;
    _T_2696_im <= _T_2695_im;
    _T_2697_re <= _T_2696_re;
    _T_2697_im <= _T_2696_im;
    _T_2698_re <= _T_2697_re;
    _T_2698_im <= _T_2697_im;
    _T_2699_re <= _T_2698_re;
    _T_2699_im <= _T_2698_im;
    _T_2700_re <= _T_2699_re;
    _T_2700_im <= _T_2699_im;
    _T_2701_re <= _T_2700_re;
    _T_2701_im <= _T_2700_im;
    _T_2702_re <= _T_2701_re;
    _T_2702_im <= _T_2701_im;
    _T_2703_re <= _T_2702_re;
    _T_2703_im <= _T_2702_im;
    _T_2704_re <= _T_2703_re;
    _T_2704_im <= _T_2703_im;
    _T_2705_re <= _T_2704_re;
    _T_2705_im <= _T_2704_im;
    _T_2706_re <= _T_2705_re;
    _T_2706_im <= _T_2705_im;
    _T_2707_re <= _T_2706_re;
    _T_2707_im <= _T_2706_im;
    _T_2708_re <= _T_2707_re;
    _T_2708_im <= _T_2707_im;
    _T_2709_re <= _T_2708_re;
    _T_2709_im <= _T_2708_im;
    _T_2710_re <= _T_2709_re;
    _T_2710_im <= _T_2709_im;
    _T_2711_re <= _T_2710_re;
    _T_2711_im <= _T_2710_im;
    _T_2712_re <= _T_2711_re;
    _T_2712_im <= _T_2711_im;
    _T_2713_re <= _T_2712_re;
    _T_2713_im <= _T_2712_im;
    _T_2714_re <= _T_2713_re;
    _T_2714_im <= _T_2713_im;
    _T_2715_re <= _T_2714_re;
    _T_2715_im <= _T_2714_im;
    _T_2716_re <= _T_2715_re;
    _T_2716_im <= _T_2715_im;
    _T_2717_re <= _T_2716_re;
    _T_2717_im <= _T_2716_im;
    _T_2718_re <= _T_2717_re;
    _T_2718_im <= _T_2717_im;
    _T_2719_re <= _T_2718_re;
    _T_2719_im <= _T_2718_im;
    _T_2720_re <= _T_2719_re;
    _T_2720_im <= _T_2719_im;
    _T_2721_re <= _T_2720_re;
    _T_2721_im <= _T_2720_im;
    _T_2722_re <= _T_2721_re;
    _T_2722_im <= _T_2721_im;
    _T_2723_re <= _T_2722_re;
    _T_2723_im <= _T_2722_im;
    _T_2724_re <= _T_2723_re;
    _T_2724_im <= _T_2723_im;
    _T_2725_re <= _T_2724_re;
    _T_2725_im <= _T_2724_im;
    _T_2726_re <= _T_2725_re;
    _T_2726_im <= _T_2725_im;
    _T_2727_re <= _T_2726_re;
    _T_2727_im <= _T_2726_im;
    _T_2728_re <= _T_2727_re;
    _T_2728_im <= _T_2727_im;
    _T_2729_re <= _T_2728_re;
    _T_2729_im <= _T_2728_im;
    _T_2730_re <= _T_2729_re;
    _T_2730_im <= _T_2729_im;
    _T_2731_re <= _T_2730_re;
    _T_2731_im <= _T_2730_im;
    _T_2732_re <= _T_2731_re;
    _T_2732_im <= _T_2731_im;
    _T_2733_re <= _T_2732_re;
    _T_2733_im <= _T_2732_im;
    _T_2734_re <= _T_2733_re;
    _T_2734_im <= _T_2733_im;
    _T_2735_re <= _T_2734_re;
    _T_2735_im <= _T_2734_im;
    _T_2736_re <= _T_2735_re;
    _T_2736_im <= _T_2735_im;
    _T_2737_re <= _T_2736_re;
    _T_2737_im <= _T_2736_im;
    _T_2738_re <= _T_2737_re;
    _T_2738_im <= _T_2737_im;
    _T_2739_re <= _T_2738_re;
    _T_2739_im <= _T_2738_im;
    _T_2740_re <= _T_2739_re;
    _T_2740_im <= _T_2739_im;
    _T_2741_re <= _T_2740_re;
    _T_2741_im <= _T_2740_im;
    _T_2742_re <= _T_2741_re;
    _T_2742_im <= _T_2741_im;
    _T_2743_re <= _T_2742_re;
    _T_2743_im <= _T_2742_im;
    _T_2744_re <= _T_2743_re;
    _T_2744_im <= _T_2743_im;
    _T_2745_re <= _T_2744_re;
    _T_2745_im <= _T_2744_im;
    _T_2746_re <= _T_2745_re;
    _T_2746_im <= _T_2745_im;
    _T_2747_re <= _T_2746_re;
    _T_2747_im <= _T_2746_im;
    _T_2748_re <= _T_2747_re;
    _T_2748_im <= _T_2747_im;
    _T_2749_re <= _T_2748_re;
    _T_2749_im <= _T_2748_im;
    _T_2750_re <= _T_2749_re;
    _T_2750_im <= _T_2749_im;
    _T_2751_re <= _T_2750_re;
    _T_2751_im <= _T_2750_im;
    _T_2752_re <= _T_2751_re;
    _T_2752_im <= _T_2751_im;
    _T_2753_re <= _T_2752_re;
    _T_2753_im <= _T_2752_im;
    _T_2754_re <= _T_2753_re;
    _T_2754_im <= _T_2753_im;
    _T_2755_re <= _T_2754_re;
    _T_2755_im <= _T_2754_im;
    _T_2756_re <= _T_2755_re;
    _T_2756_im <= _T_2755_im;
    _T_2757_re <= _T_2756_re;
    _T_2757_im <= _T_2756_im;
    _T_2758_re <= _T_2757_re;
    _T_2758_im <= _T_2757_im;
    _T_2759_re <= _T_2758_re;
    _T_2759_im <= _T_2758_im;
    _T_2760_re <= _T_2759_re;
    _T_2760_im <= _T_2759_im;
    _T_2761_re <= _T_2760_re;
    _T_2761_im <= _T_2760_im;
    _T_2762_re <= _T_2761_re;
    _T_2762_im <= _T_2761_im;
    _T_2763_re <= _T_2762_re;
    _T_2763_im <= _T_2762_im;
    _T_2764_re <= _T_2763_re;
    _T_2764_im <= _T_2763_im;
    _T_2765_re <= _T_2764_re;
    _T_2765_im <= _T_2764_im;
    _T_2766_re <= _T_2765_re;
    _T_2766_im <= _T_2765_im;
    _T_2767_re <= _T_2766_re;
    _T_2767_im <= _T_2766_im;
    _T_2768_re <= _T_2767_re;
    _T_2768_im <= _T_2767_im;
    _T_2769_re <= _T_2768_re;
    _T_2769_im <= _T_2768_im;
    _T_2770_re <= _T_2769_re;
    _T_2770_im <= _T_2769_im;
    _T_2771_re <= _T_2770_re;
    _T_2771_im <= _T_2770_im;
    _T_2772_re <= _T_2771_re;
    _T_2772_im <= _T_2771_im;
    _T_2773_re <= _T_2772_re;
    _T_2773_im <= _T_2772_im;
    _T_2774_re <= _T_2773_re;
    _T_2774_im <= _T_2773_im;
    _T_2775_re <= _T_2774_re;
    _T_2775_im <= _T_2774_im;
    _T_2776_re <= _T_2775_re;
    _T_2776_im <= _T_2775_im;
    _T_2777_re <= _T_2776_re;
    _T_2777_im <= _T_2776_im;
    _T_2778_re <= _T_2777_re;
    _T_2778_im <= _T_2777_im;
    _T_2779_re <= _T_2778_re;
    _T_2779_im <= _T_2778_im;
    _T_2780_re <= _T_2779_re;
    _T_2780_im <= _T_2779_im;
    _T_2781_re <= _T_2780_re;
    _T_2781_im <= _T_2780_im;
    _T_2782_re <= _T_2781_re;
    _T_2782_im <= _T_2781_im;
    _T_2783_re <= _T_2782_re;
    _T_2783_im <= _T_2782_im;
    _T_2784_re <= _T_2783_re;
    _T_2784_im <= _T_2783_im;
    _T_2785_re <= _T_2784_re;
    _T_2785_im <= _T_2784_im;
    _T_2786_re <= _T_2785_re;
    _T_2786_im <= _T_2785_im;
    _T_2787_re <= _T_2786_re;
    _T_2787_im <= _T_2786_im;
    _T_2788_re <= _T_2787_re;
    _T_2788_im <= _T_2787_im;
    _T_2789_re <= _T_2788_re;
    _T_2789_im <= _T_2788_im;
    _T_2790_re <= _T_2789_re;
    _T_2790_im <= _T_2789_im;
    _T_2791_re <= _T_2790_re;
    _T_2791_im <= _T_2790_im;
    _T_2792_re <= _T_2791_re;
    _T_2792_im <= _T_2791_im;
    _T_2793_re <= _T_2792_re;
    _T_2793_im <= _T_2792_im;
    _T_2794_re <= _T_2793_re;
    _T_2794_im <= _T_2793_im;
    _T_2795_re <= _T_2794_re;
    _T_2795_im <= _T_2794_im;
    _T_2796_re <= _T_2795_re;
    _T_2796_im <= _T_2795_im;
    _T_2797_re <= _T_2796_re;
    _T_2797_im <= _T_2796_im;
    _T_2798_re <= _T_2797_re;
    _T_2798_im <= _T_2797_im;
    _T_2799_re <= _T_2798_re;
    _T_2799_im <= _T_2798_im;
    _T_2800_re <= _T_2799_re;
    _T_2800_im <= _T_2799_im;
    _T_2801_re <= _T_2800_re;
    _T_2801_im <= _T_2800_im;
    _T_2802_re <= _T_2801_re;
    _T_2802_im <= _T_2801_im;
    _T_2803_re <= _T_2802_re;
    _T_2803_im <= _T_2802_im;
    _T_2804_re <= _T_2803_re;
    _T_2804_im <= _T_2803_im;
    _T_2805_re <= _T_2804_re;
    _T_2805_im <= _T_2804_im;
    _T_2806_re <= _T_2805_re;
    _T_2806_im <= _T_2805_im;
    _T_2807_re <= _T_2806_re;
    _T_2807_im <= _T_2806_im;
    _T_2808_re <= _T_2807_re;
    _T_2808_im <= _T_2807_im;
    _T_2809_re <= _T_2808_re;
    _T_2809_im <= _T_2808_im;
    _T_2810_re <= _T_2809_re;
    _T_2810_im <= _T_2809_im;
    _T_2811_re <= _T_2810_re;
    _T_2811_im <= _T_2810_im;
    _T_2812_re <= _T_2811_re;
    _T_2812_im <= _T_2811_im;
    _T_2813_re <= _T_2812_re;
    _T_2813_im <= _T_2812_im;
    _T_2814_re <= _T_2813_re;
    _T_2814_im <= _T_2813_im;
    _T_2815_re <= _T_2814_re;
    _T_2815_im <= _T_2814_im;
    _T_2816_re <= _T_2815_re;
    _T_2816_im <= _T_2815_im;
    _T_2817_re <= _T_2816_re;
    _T_2817_im <= _T_2816_im;
    _T_2818_re <= _T_2817_re;
    _T_2818_im <= _T_2817_im;
    _T_2819_re <= _T_2818_re;
    _T_2819_im <= _T_2818_im;
    _T_2820_re <= _T_2819_re;
    _T_2820_im <= _T_2819_im;
    _T_2821_re <= _T_2820_re;
    _T_2821_im <= _T_2820_im;
    _T_2822_re <= _T_2821_re;
    _T_2822_im <= _T_2821_im;
    _T_2823_re <= _T_2822_re;
    _T_2823_im <= _T_2822_im;
    _T_2824_re <= _T_2823_re;
    _T_2824_im <= _T_2823_im;
    _T_2825_re <= _T_2824_re;
    _T_2825_im <= _T_2824_im;
    _T_2826_re <= _T_2825_re;
    _T_2826_im <= _T_2825_im;
    _T_2827_re <= _T_2826_re;
    _T_2827_im <= _T_2826_im;
    _T_2828_re <= _T_2827_re;
    _T_2828_im <= _T_2827_im;
    _T_2829_re <= _T_2828_re;
    _T_2829_im <= _T_2828_im;
    _T_2830_re <= _T_2829_re;
    _T_2830_im <= _T_2829_im;
    _T_2831_re <= _T_2830_re;
    _T_2831_im <= _T_2830_im;
    _T_2832_re <= _T_2831_re;
    _T_2832_im <= _T_2831_im;
    _T_2833_re <= _T_2832_re;
    _T_2833_im <= _T_2832_im;
    _T_2834_re <= _T_2833_re;
    _T_2834_im <= _T_2833_im;
    _T_2835_re <= _T_2834_re;
    _T_2835_im <= _T_2834_im;
    _T_2836_re <= _T_2835_re;
    _T_2836_im <= _T_2835_im;
    _T_2837_re <= _T_2836_re;
    _T_2837_im <= _T_2836_im;
    _T_2838_re <= _T_2837_re;
    _T_2838_im <= _T_2837_im;
    _T_2839_re <= _T_2838_re;
    _T_2839_im <= _T_2838_im;
    _T_2840_re <= _T_2839_re;
    _T_2840_im <= _T_2839_im;
    _T_2841_re <= _T_2840_re;
    _T_2841_im <= _T_2840_im;
    _T_2842_re <= _T_2841_re;
    _T_2842_im <= _T_2841_im;
    _T_2843_re <= _T_2842_re;
    _T_2843_im <= _T_2842_im;
    _T_2844_re <= _T_2843_re;
    _T_2844_im <= _T_2843_im;
    _T_2845_re <= _T_2844_re;
    _T_2845_im <= _T_2844_im;
    _T_2846_re <= _T_2845_re;
    _T_2846_im <= _T_2845_im;
    _T_2847_re <= _T_2846_re;
    _T_2847_im <= _T_2846_im;
    _T_2848_re <= _T_2847_re;
    _T_2848_im <= _T_2847_im;
    _T_2849_re <= _T_2848_re;
    _T_2849_im <= _T_2848_im;
    _T_2850_re <= _T_2849_re;
    _T_2850_im <= _T_2849_im;
    _T_2851_re <= _T_2850_re;
    _T_2851_im <= _T_2850_im;
    _T_2852_re <= _T_2851_re;
    _T_2852_im <= _T_2851_im;
    _T_2853_re <= _T_2852_re;
    _T_2853_im <= _T_2852_im;
    _T_2854_re <= _T_2853_re;
    _T_2854_im <= _T_2853_im;
    _T_2855_re <= _T_2854_re;
    _T_2855_im <= _T_2854_im;
    _T_2856_re <= _T_2855_re;
    _T_2856_im <= _T_2855_im;
    _T_2857_re <= _T_2856_re;
    _T_2857_im <= _T_2856_im;
    _T_2858_re <= _T_2857_re;
    _T_2858_im <= _T_2857_im;
    _T_2859_re <= _T_2858_re;
    _T_2859_im <= _T_2858_im;
    _T_2860_re <= _T_2859_re;
    _T_2860_im <= _T_2859_im;
    _T_2861_re <= _T_2860_re;
    _T_2861_im <= _T_2860_im;
    _T_2862_re <= _T_2861_re;
    _T_2862_im <= _T_2861_im;
    _T_2863_re <= _T_2862_re;
    _T_2863_im <= _T_2862_im;
    _T_2864_re <= _T_2863_re;
    _T_2864_im <= _T_2863_im;
    _T_2865_re <= _T_2864_re;
    _T_2865_im <= _T_2864_im;
    _T_2866_re <= _T_2865_re;
    _T_2866_im <= _T_2865_im;
    _T_2867_re <= _T_2866_re;
    _T_2867_im <= _T_2866_im;
    _T_2868_re <= _T_2867_re;
    _T_2868_im <= _T_2867_im;
    _T_2869_re <= _T_2868_re;
    _T_2869_im <= _T_2868_im;
    _T_2870_re <= _T_2869_re;
    _T_2870_im <= _T_2869_im;
    _T_2871_re <= _T_2870_re;
    _T_2871_im <= _T_2870_im;
    _T_2872_re <= _T_2871_re;
    _T_2872_im <= _T_2871_im;
    _T_2873_re <= _T_2872_re;
    _T_2873_im <= _T_2872_im;
    _T_2874_re <= _T_2873_re;
    _T_2874_im <= _T_2873_im;
    _T_2875_re <= _T_2874_re;
    _T_2875_im <= _T_2874_im;
    _T_2876_re <= _T_2875_re;
    _T_2876_im <= _T_2875_im;
    _T_2877_re <= _T_2876_re;
    _T_2877_im <= _T_2876_im;
    _T_2878_re <= _T_2877_re;
    _T_2878_im <= _T_2877_im;
    _T_2879_re <= _T_2878_re;
    _T_2879_im <= _T_2878_im;
    _T_2880_re <= _T_2879_re;
    _T_2880_im <= _T_2879_im;
    _T_2881_re <= _T_2880_re;
    _T_2881_im <= _T_2880_im;
    _T_2882_re <= _T_2881_re;
    _T_2882_im <= _T_2881_im;
    _T_2883_re <= _T_2882_re;
    _T_2883_im <= _T_2882_im;
    _T_2884_re <= _T_2883_re;
    _T_2884_im <= _T_2883_im;
    _T_2885_re <= _T_2884_re;
    _T_2885_im <= _T_2884_im;
    _T_2886_re <= _T_2885_re;
    _T_2886_im <= _T_2885_im;
    _T_2887_re <= _T_2886_re;
    _T_2887_im <= _T_2886_im;
    _T_2888_re <= _T_2887_re;
    _T_2888_im <= _T_2887_im;
    _T_2889_re <= _T_2888_re;
    _T_2889_im <= _T_2888_im;
    _T_2890_re <= _T_2889_re;
    _T_2890_im <= _T_2889_im;
    _T_2891_re <= _T_2890_re;
    _T_2891_im <= _T_2890_im;
    _T_2892_re <= _T_2891_re;
    _T_2892_im <= _T_2891_im;
    _T_2893_re <= _T_2892_re;
    _T_2893_im <= _T_2892_im;
    _T_2894_re <= _T_2893_re;
    _T_2894_im <= _T_2893_im;
    _T_2895_re <= _T_2894_re;
    _T_2895_im <= _T_2894_im;
    _T_2896_re <= _T_2895_re;
    _T_2896_im <= _T_2895_im;
    _T_2897_re <= _T_2896_re;
    _T_2897_im <= _T_2896_im;
    _T_2898_re <= _T_2897_re;
    _T_2898_im <= _T_2897_im;
    _T_2899_re <= _T_2898_re;
    _T_2899_im <= _T_2898_im;
    _T_2900_re <= _T_2899_re;
    _T_2900_im <= _T_2899_im;
    _T_2901_re <= _T_2900_re;
    _T_2901_im <= _T_2900_im;
    _T_2902_re <= _T_2901_re;
    _T_2902_im <= _T_2901_im;
    _T_2903_re <= _T_2902_re;
    _T_2903_im <= _T_2902_im;
    _T_2904_re <= _T_2903_re;
    _T_2904_im <= _T_2903_im;
    _T_2905_re <= _T_2904_re;
    _T_2905_im <= _T_2904_im;
    _T_2906_re <= _T_2905_re;
    _T_2906_im <= _T_2905_im;
    _T_2907_re <= _T_2906_re;
    _T_2907_im <= _T_2906_im;
    _T_2908_re <= _T_2907_re;
    _T_2908_im <= _T_2907_im;
    _T_2909_re <= _T_2908_re;
    _T_2909_im <= _T_2908_im;
    _T_2910_re <= _T_2909_re;
    _T_2910_im <= _T_2909_im;
    _T_2911_re <= _T_2910_re;
    _T_2911_im <= _T_2910_im;
    _T_2912_re <= _T_2911_re;
    _T_2912_im <= _T_2911_im;
    _T_2913_re <= _T_2912_re;
    _T_2913_im <= _T_2912_im;
    _T_2914_re <= _T_2913_re;
    _T_2914_im <= _T_2913_im;
    _T_2915_re <= _T_2914_re;
    _T_2915_im <= _T_2914_im;
    _T_2916_re <= _T_2915_re;
    _T_2916_im <= _T_2915_im;
    _T_2917_re <= _T_2916_re;
    _T_2917_im <= _T_2916_im;
    _T_2918_re <= _T_2917_re;
    _T_2918_im <= _T_2917_im;
    _T_2919_re <= _T_2918_re;
    _T_2919_im <= _T_2918_im;
    _T_2920_re <= _T_2919_re;
    _T_2920_im <= _T_2919_im;
    _T_2921_re <= _T_2920_re;
    _T_2921_im <= _T_2920_im;
    _T_2922_re <= _T_2921_re;
    _T_2922_im <= _T_2921_im;
    _T_2923_re <= _T_2922_re;
    _T_2923_im <= _T_2922_im;
    _T_2924_re <= _T_2923_re;
    _T_2924_im <= _T_2923_im;
    _T_2925_re <= _T_2924_re;
    _T_2925_im <= _T_2924_im;
    _T_2926_re <= _T_2925_re;
    _T_2926_im <= _T_2925_im;
    _T_2927_re <= _T_2926_re;
    _T_2927_im <= _T_2926_im;
    _T_2928_re <= _T_2927_re;
    _T_2928_im <= _T_2927_im;
    _T_2929_re <= _T_2928_re;
    _T_2929_im <= _T_2928_im;
    _T_2930_re <= _T_2929_re;
    _T_2930_im <= _T_2929_im;
    _T_2931_re <= _T_2930_re;
    _T_2931_im <= _T_2930_im;
    _T_2932_re <= _T_2931_re;
    _T_2932_im <= _T_2931_im;
    _T_2933_re <= _T_2932_re;
    _T_2933_im <= _T_2932_im;
    _T_2934_re <= _T_2933_re;
    _T_2934_im <= _T_2933_im;
    _T_2935_re <= _T_2934_re;
    _T_2935_im <= _T_2934_im;
    _T_2936_re <= _T_2935_re;
    _T_2936_im <= _T_2935_im;
    _T_2937_re <= _T_2936_re;
    _T_2937_im <= _T_2936_im;
    _T_2938_re <= _T_2937_re;
    _T_2938_im <= _T_2937_im;
    _T_2939_re <= _T_2938_re;
    _T_2939_im <= _T_2938_im;
    _T_2940_re <= _T_2939_re;
    _T_2940_im <= _T_2939_im;
    _T_2941_re <= _T_2940_re;
    _T_2941_im <= _T_2940_im;
    _T_2942_re <= _T_2941_re;
    _T_2942_im <= _T_2941_im;
    _T_2943_re <= _T_2942_re;
    _T_2943_im <= _T_2942_im;
    _T_2944_re <= _T_2943_re;
    _T_2944_im <= _T_2943_im;
    _T_2945_re <= _T_2944_re;
    _T_2945_im <= _T_2944_im;
    _T_2946_re <= _T_2945_re;
    _T_2946_im <= _T_2945_im;
    _T_2947_re <= _T_2946_re;
    _T_2947_im <= _T_2946_im;
    _T_2948_re <= _T_2947_re;
    _T_2948_im <= _T_2947_im;
    _T_2949_re <= _T_2948_re;
    _T_2949_im <= _T_2948_im;
    _T_2950_re <= _T_2949_re;
    _T_2950_im <= _T_2949_im;
    _T_2951_re <= _T_2950_re;
    _T_2951_im <= _T_2950_im;
    _T_2952_re <= _T_2951_re;
    _T_2952_im <= _T_2951_im;
    _T_2953_re <= _T_2952_re;
    _T_2953_im <= _T_2952_im;
    _T_2954_re <= _T_2953_re;
    _T_2954_im <= _T_2953_im;
    _T_2955_re <= _T_2954_re;
    _T_2955_im <= _T_2954_im;
    _T_2956_re <= _T_2955_re;
    _T_2956_im <= _T_2955_im;
    _T_2957_re <= _T_2956_re;
    _T_2957_im <= _T_2956_im;
    _T_2958_re <= _T_2957_re;
    _T_2958_im <= _T_2957_im;
    _T_2959_re <= _T_2958_re;
    _T_2959_im <= _T_2958_im;
    _T_2960_re <= _T_2959_re;
    _T_2960_im <= _T_2959_im;
    _T_2961_re <= _T_2960_re;
    _T_2961_im <= _T_2960_im;
    _T_2962_re <= _T_2961_re;
    _T_2962_im <= _T_2961_im;
    _T_2963_re <= _T_2962_re;
    _T_2963_im <= _T_2962_im;
    _T_2964_re <= _T_2963_re;
    _T_2964_im <= _T_2963_im;
    _T_2965_re <= _T_2964_re;
    _T_2965_im <= _T_2964_im;
    _T_2966_re <= _T_2965_re;
    _T_2966_im <= _T_2965_im;
    _T_2967_re <= _T_2966_re;
    _T_2967_im <= _T_2966_im;
    _T_2968_re <= _T_2967_re;
    _T_2968_im <= _T_2967_im;
    _T_2969_re <= _T_2968_re;
    _T_2969_im <= _T_2968_im;
    _T_2970_re <= _T_2969_re;
    _T_2970_im <= _T_2969_im;
    _T_2971_re <= _T_2970_re;
    _T_2971_im <= _T_2970_im;
    _T_2972_re <= _T_2971_re;
    _T_2972_im <= _T_2971_im;
    _T_2973_re <= _T_2972_re;
    _T_2973_im <= _T_2972_im;
    _T_2974_re <= _T_2973_re;
    _T_2974_im <= _T_2973_im;
    _T_2975_re <= _T_2974_re;
    _T_2975_im <= _T_2974_im;
    _T_2976_re <= _T_2975_re;
    _T_2976_im <= _T_2975_im;
    _T_2977_re <= _T_2976_re;
    _T_2977_im <= _T_2976_im;
    _T_2978_re <= _T_2977_re;
    _T_2978_im <= _T_2977_im;
    _T_2979_re <= _T_2978_re;
    _T_2979_im <= _T_2978_im;
    _T_2980_re <= _T_2979_re;
    _T_2980_im <= _T_2979_im;
    _T_2981_re <= _T_2980_re;
    _T_2981_im <= _T_2980_im;
    _T_2982_re <= _T_2981_re;
    _T_2982_im <= _T_2981_im;
    _T_2983_re <= _T_2982_re;
    _T_2983_im <= _T_2982_im;
    _T_2984_re <= _T_2983_re;
    _T_2984_im <= _T_2983_im;
    _T_2985_re <= _T_2984_re;
    _T_2985_im <= _T_2984_im;
    _T_2986_re <= _T_2985_re;
    _T_2986_im <= _T_2985_im;
    _T_2987_re <= _T_2986_re;
    _T_2987_im <= _T_2986_im;
    _T_2988_re <= _T_2987_re;
    _T_2988_im <= _T_2987_im;
    _T_2989_re <= _T_2988_re;
    _T_2989_im <= _T_2988_im;
    _T_2990_re <= _T_2989_re;
    _T_2990_im <= _T_2989_im;
    _T_2991_re <= _T_2990_re;
    _T_2991_im <= _T_2990_im;
    _T_2992_re <= _T_2991_re;
    _T_2992_im <= _T_2991_im;
    _T_2993_re <= _T_2992_re;
    _T_2993_im <= _T_2992_im;
    _T_2994_re <= _T_2993_re;
    _T_2994_im <= _T_2993_im;
    _T_2995_re <= _T_2994_re;
    _T_2995_im <= _T_2994_im;
    _T_2996_re <= _T_2995_re;
    _T_2996_im <= _T_2995_im;
    _T_2997_re <= _T_2996_re;
    _T_2997_im <= _T_2996_im;
    _T_2998_re <= _T_2997_re;
    _T_2998_im <= _T_2997_im;
    _T_2999_re <= _T_2998_re;
    _T_2999_im <= _T_2998_im;
    _T_3000_re <= _T_2999_re;
    _T_3000_im <= _T_2999_im;
    _T_3001_re <= _T_3000_re;
    _T_3001_im <= _T_3000_im;
    _T_3002_re <= _T_3001_re;
    _T_3002_im <= _T_3001_im;
    _T_3003_re <= _T_3002_re;
    _T_3003_im <= _T_3002_im;
    _T_3004_re <= _T_3003_re;
    _T_3004_im <= _T_3003_im;
    _T_3005_re <= _T_3004_re;
    _T_3005_im <= _T_3004_im;
    _T_3006_re <= _T_3005_re;
    _T_3006_im <= _T_3005_im;
    _T_3007_re <= _T_3006_re;
    _T_3007_im <= _T_3006_im;
    _T_3008_re <= _T_3007_re;
    _T_3008_im <= _T_3007_im;
    _T_3009_re <= _T_3008_re;
    _T_3009_im <= _T_3008_im;
    _T_3010_re <= _T_3009_re;
    _T_3010_im <= _T_3009_im;
    _T_3011_re <= _T_3010_re;
    _T_3011_im <= _T_3010_im;
    _T_3012_re <= _T_3011_re;
    _T_3012_im <= _T_3011_im;
    _T_3013_re <= _T_3012_re;
    _T_3013_im <= _T_3012_im;
    _T_3014_re <= _T_3013_re;
    _T_3014_im <= _T_3013_im;
    _T_3015_re <= _T_3014_re;
    _T_3015_im <= _T_3014_im;
    _T_3016_re <= _T_3015_re;
    _T_3016_im <= _T_3015_im;
    _T_3017_re <= _T_3016_re;
    _T_3017_im <= _T_3016_im;
    _T_3018_re <= _T_3017_re;
    _T_3018_im <= _T_3017_im;
    _T_3019_re <= _T_3018_re;
    _T_3019_im <= _T_3018_im;
    _T_3020_re <= _T_3019_re;
    _T_3020_im <= _T_3019_im;
    _T_3021_re <= _T_3020_re;
    _T_3021_im <= _T_3020_im;
    _T_3022_re <= _T_3021_re;
    _T_3022_im <= _T_3021_im;
    _T_3023_re <= _T_3022_re;
    _T_3023_im <= _T_3022_im;
    _T_3024_re <= _T_3023_re;
    _T_3024_im <= _T_3023_im;
    _T_3025_re <= _T_3024_re;
    _T_3025_im <= _T_3024_im;
    _T_3026_re <= _T_3025_re;
    _T_3026_im <= _T_3025_im;
    _T_3027_re <= _T_3026_re;
    _T_3027_im <= _T_3026_im;
    _T_3028_re <= _T_3027_re;
    _T_3028_im <= _T_3027_im;
    _T_3029_re <= _T_3028_re;
    _T_3029_im <= _T_3028_im;
    _T_3030_re <= _T_3029_re;
    _T_3030_im <= _T_3029_im;
    _T_3031_re <= _T_3030_re;
    _T_3031_im <= _T_3030_im;
    _T_3032_re <= _T_3031_re;
    _T_3032_im <= _T_3031_im;
    _T_3033_re <= _T_3032_re;
    _T_3033_im <= _T_3032_im;
    _T_3034_re <= _T_3033_re;
    _T_3034_im <= _T_3033_im;
    _T_3035_re <= _T_3034_re;
    _T_3035_im <= _T_3034_im;
    _T_3036_re <= _T_3035_re;
    _T_3036_im <= _T_3035_im;
    _T_3037_re <= _T_3036_re;
    _T_3037_im <= _T_3036_im;
    _T_3038_re <= _T_3037_re;
    _T_3038_im <= _T_3037_im;
    _T_3039_re <= _T_3038_re;
    _T_3039_im <= _T_3038_im;
    _T_3040_re <= _T_3039_re;
    _T_3040_im <= _T_3039_im;
    _T_3041_re <= _T_3040_re;
    _T_3041_im <= _T_3040_im;
    _T_3042_re <= _T_3041_re;
    _T_3042_im <= _T_3041_im;
    _T_3043_re <= _T_3042_re;
    _T_3043_im <= _T_3042_im;
    _T_3044_re <= _T_3043_re;
    _T_3044_im <= _T_3043_im;
    _T_3045_re <= _T_3044_re;
    _T_3045_im <= _T_3044_im;
    _T_3046_re <= _T_3045_re;
    _T_3046_im <= _T_3045_im;
    _T_3047_re <= _T_3046_re;
    _T_3047_im <= _T_3046_im;
    _T_3048_re <= _T_3047_re;
    _T_3048_im <= _T_3047_im;
    _T_3049_re <= _T_3048_re;
    _T_3049_im <= _T_3048_im;
    _T_3050_re <= _T_3049_re;
    _T_3050_im <= _T_3049_im;
    _T_3051_re <= _T_3050_re;
    _T_3051_im <= _T_3050_im;
    _T_3052_re <= _T_3051_re;
    _T_3052_im <= _T_3051_im;
    _T_3053_re <= _T_3052_re;
    _T_3053_im <= _T_3052_im;
    _T_3054_re <= _T_3053_re;
    _T_3054_im <= _T_3053_im;
    _T_3055_re <= _T_3054_re;
    _T_3055_im <= _T_3054_im;
    _T_3056_re <= _T_3055_re;
    _T_3056_im <= _T_3055_im;
    _T_3057_re <= _T_3056_re;
    _T_3057_im <= _T_3056_im;
    _T_3058_re <= _T_3057_re;
    _T_3058_im <= _T_3057_im;
    _T_3059_re <= _T_3058_re;
    _T_3059_im <= _T_3058_im;
    _T_3060_re <= _T_3059_re;
    _T_3060_im <= _T_3059_im;
    _T_3061_re <= _T_3060_re;
    _T_3061_im <= _T_3060_im;
    _T_3062_re <= _T_3061_re;
    _T_3062_im <= _T_3061_im;
    _T_3063_re <= _T_3062_re;
    _T_3063_im <= _T_3062_im;
    _T_3064_re <= _T_3063_re;
    _T_3064_im <= _T_3063_im;
    _T_3065_re <= _T_3064_re;
    _T_3065_im <= _T_3064_im;
    _T_3066_re <= _T_3065_re;
    _T_3066_im <= _T_3065_im;
    _T_3067_re <= _T_3066_re;
    _T_3067_im <= _T_3066_im;
    _T_3068_re <= _T_3067_re;
    _T_3068_im <= _T_3067_im;
    _T_3069_re <= _T_3068_re;
    _T_3069_im <= _T_3068_im;
    _T_3070_re <= _T_3069_re;
    _T_3070_im <= _T_3069_im;
    _T_3071_re <= _T_3070_re;
    _T_3071_im <= _T_3070_im;
    _T_3072_re <= _T_3071_re;
    _T_3072_im <= _T_3071_im;
    _T_3073_re <= _T_3072_re;
    _T_3073_im <= _T_3072_im;
    _T_3074_re <= _T_3073_re;
    _T_3074_im <= _T_3073_im;
    _T_3075_re <= _T_3074_re;
    _T_3075_im <= _T_3074_im;
    _T_3076_re <= _T_3075_re;
    _T_3076_im <= _T_3075_im;
    _T_3077_re <= _T_3076_re;
    _T_3077_im <= _T_3076_im;
    _T_3078_re <= _T_3077_re;
    _T_3078_im <= _T_3077_im;
    _T_3079_re <= _T_3078_re;
    _T_3079_im <= _T_3078_im;
    _T_3080_re <= _T_3079_re;
    _T_3080_im <= _T_3079_im;
    _T_3081_re <= _T_3080_re;
    _T_3081_im <= _T_3080_im;
    _T_3082_re <= _T_3081_re;
    _T_3082_im <= _T_3081_im;
    _T_3083_re <= _T_3082_re;
    _T_3083_im <= _T_3082_im;
    _T_3084_re <= _T_3083_re;
    _T_3084_im <= _T_3083_im;
    _T_3085_re <= _T_3084_re;
    _T_3085_im <= _T_3084_im;
    _T_3086_re <= _T_3085_re;
    _T_3086_im <= _T_3085_im;
    _T_3087_re <= _T_3086_re;
    _T_3087_im <= _T_3086_im;
    _T_3088_re <= _T_3087_re;
    _T_3088_im <= _T_3087_im;
    _T_3089_re <= _T_3088_re;
    _T_3089_im <= _T_3088_im;
    _T_3090_re <= _T_3089_re;
    _T_3090_im <= _T_3089_im;
    _T_3091_re <= _T_3090_re;
    _T_3091_im <= _T_3090_im;
    _T_3092_re <= _T_3091_re;
    _T_3092_im <= _T_3091_im;
    _T_3093_re <= _T_3092_re;
    _T_3093_im <= _T_3092_im;
    _T_3094_re <= _T_3093_re;
    _T_3094_im <= _T_3093_im;
    _T_3095_re <= _T_3094_re;
    _T_3095_im <= _T_3094_im;
    _T_3096_re <= _T_3095_re;
    _T_3096_im <= _T_3095_im;
    _T_3097_re <= _T_3096_re;
    _T_3097_im <= _T_3096_im;
    _T_3098_re <= _T_3097_re;
    _T_3098_im <= _T_3097_im;
    _T_3099_re <= _T_3098_re;
    _T_3099_im <= _T_3098_im;
    _T_3100_re <= _T_3099_re;
    _T_3100_im <= _T_3099_im;
    _T_3101_re <= _T_3100_re;
    _T_3101_im <= _T_3100_im;
    _T_3102_re <= _T_3101_re;
    _T_3102_im <= _T_3101_im;
    _T_3103_re <= _T_3102_re;
    _T_3103_im <= _T_3102_im;
    _T_3104_re <= _T_3103_re;
    _T_3104_im <= _T_3103_im;
    _T_3105_re <= _T_3104_re;
    _T_3105_im <= _T_3104_im;
    _T_3106_re <= _T_3105_re;
    _T_3106_im <= _T_3105_im;
    _T_3107_re <= _T_3106_re;
    _T_3107_im <= _T_3106_im;
    _T_3108_re <= _T_3107_re;
    _T_3108_im <= _T_3107_im;
    _T_3109_re <= _T_3108_re;
    _T_3109_im <= _T_3108_im;
    _T_3110_re <= _T_3109_re;
    _T_3110_im <= _T_3109_im;
    _T_3111_re <= _T_3110_re;
    _T_3111_im <= _T_3110_im;
    _T_3112_re <= _T_3111_re;
    _T_3112_im <= _T_3111_im;
    _T_3113_re <= _T_3112_re;
    _T_3113_im <= _T_3112_im;
    _T_3114_re <= _T_3113_re;
    _T_3114_im <= _T_3113_im;
    _T_3115_re <= _T_3114_re;
    _T_3115_im <= _T_3114_im;
    _T_3116_re <= _T_3115_re;
    _T_3116_im <= _T_3115_im;
    _T_3117_re <= _T_3116_re;
    _T_3117_im <= _T_3116_im;
    _T_3118_re <= _T_3117_re;
    _T_3118_im <= _T_3117_im;
    _T_3119_re <= _T_3118_re;
    _T_3119_im <= _T_3118_im;
    _T_3120_re <= _T_3119_re;
    _T_3120_im <= _T_3119_im;
    _T_3121_re <= _T_3120_re;
    _T_3121_im <= _T_3120_im;
    _T_3122_re <= _T_3121_re;
    _T_3122_im <= _T_3121_im;
    _T_3123_re <= _T_3122_re;
    _T_3123_im <= _T_3122_im;
    _T_3124_re <= _T_3123_re;
    _T_3124_im <= _T_3123_im;
    _T_3125_re <= _T_3124_re;
    _T_3125_im <= _T_3124_im;
    _T_3126_re <= _T_3125_re;
    _T_3126_im <= _T_3125_im;
    _T_3127_re <= _T_3126_re;
    _T_3127_im <= _T_3126_im;
    _T_3128_re <= _T_3127_re;
    _T_3128_im <= _T_3127_im;
    _T_3129_re <= _T_3128_re;
    _T_3129_im <= _T_3128_im;
    _T_3130_re <= _T_3129_re;
    _T_3130_im <= _T_3129_im;
    _T_3131_re <= _T_3130_re;
    _T_3131_im <= _T_3130_im;
    _T_3132_re <= _T_3131_re;
    _T_3132_im <= _T_3131_im;
    _T_3133_re <= _T_3132_re;
    _T_3133_im <= _T_3132_im;
    _T_3134_re <= _T_3133_re;
    _T_3134_im <= _T_3133_im;
    _T_3135_re <= _T_3134_re;
    _T_3135_im <= _T_3134_im;
    _T_3136_re <= _T_3135_re;
    _T_3136_im <= _T_3135_im;
    _T_3137_re <= _T_3136_re;
    _T_3137_im <= _T_3136_im;
    _T_3138_re <= _T_3137_re;
    _T_3138_im <= _T_3137_im;
    _T_3139_re <= _T_3138_re;
    _T_3139_im <= _T_3138_im;
    _T_3140_re <= _T_3139_re;
    _T_3140_im <= _T_3139_im;
    _T_3141_re <= _T_3140_re;
    _T_3141_im <= _T_3140_im;
    _T_3142_re <= _T_3141_re;
    _T_3142_im <= _T_3141_im;
    _T_3143_re <= _T_3142_re;
    _T_3143_im <= _T_3142_im;
    _T_3144_re <= _T_3143_re;
    _T_3144_im <= _T_3143_im;
    _T_3145_re <= _T_3144_re;
    _T_3145_im <= _T_3144_im;
    _T_3146_re <= _T_3145_re;
    _T_3146_im <= _T_3145_im;
    _T_3147_re <= _T_3146_re;
    _T_3147_im <= _T_3146_im;
    _T_3148_re <= _T_3147_re;
    _T_3148_im <= _T_3147_im;
    _T_3149_re <= _T_3148_re;
    _T_3149_im <= _T_3148_im;
    _T_3150_re <= _T_3149_re;
    _T_3150_im <= _T_3149_im;
    _T_3151_re <= _T_3150_re;
    _T_3151_im <= _T_3150_im;
    _T_3152_re <= _T_3151_re;
    _T_3152_im <= _T_3151_im;
    _T_3153_re <= _T_3152_re;
    _T_3153_im <= _T_3152_im;
    _T_3154_re <= _T_3153_re;
    _T_3154_im <= _T_3153_im;
    _T_3155_re <= _T_3154_re;
    _T_3155_im <= _T_3154_im;
    _T_3156_re <= _T_3155_re;
    _T_3156_im <= _T_3155_im;
    _T_3157_re <= _T_3156_re;
    _T_3157_im <= _T_3156_im;
    _T_3158_re <= _T_3157_re;
    _T_3158_im <= _T_3157_im;
    _T_3159_re <= _T_3158_re;
    _T_3159_im <= _T_3158_im;
    _T_3160_re <= _T_3159_re;
    _T_3160_im <= _T_3159_im;
    _T_3161_re <= _T_3160_re;
    _T_3161_im <= _T_3160_im;
    _T_3162_re <= _T_3161_re;
    _T_3162_im <= _T_3161_im;
    _T_3163_re <= _T_3162_re;
    _T_3163_im <= _T_3162_im;
    _T_3164_re <= _T_3163_re;
    _T_3164_im <= _T_3163_im;
    _T_3165_re <= _T_3164_re;
    _T_3165_im <= _T_3164_im;
    _T_3166_re <= _T_3165_re;
    _T_3166_im <= _T_3165_im;
    _T_3167_re <= _T_3166_re;
    _T_3167_im <= _T_3166_im;
    _T_3168_re <= _T_3167_re;
    _T_3168_im <= _T_3167_im;
    _T_3169_re <= _T_3168_re;
    _T_3169_im <= _T_3168_im;
    _T_3170_re <= _T_3169_re;
    _T_3170_im <= _T_3169_im;
    _T_3171_re <= _T_3170_re;
    _T_3171_im <= _T_3170_im;
    _T_3172_re <= _T_3171_re;
    _T_3172_im <= _T_3171_im;
    _T_3173_re <= _T_3172_re;
    _T_3173_im <= _T_3172_im;
    _T_3174_re <= _T_3173_re;
    _T_3174_im <= _T_3173_im;
    _T_3175_re <= _T_3174_re;
    _T_3175_im <= _T_3174_im;
    _T_3176_re <= _T_3175_re;
    _T_3176_im <= _T_3175_im;
    _T_3177_re <= _T_3176_re;
    _T_3177_im <= _T_3176_im;
    _T_3178_re <= _T_3177_re;
    _T_3178_im <= _T_3177_im;
    _T_3179_re <= _T_3178_re;
    _T_3179_im <= _T_3178_im;
    _T_3180_re <= _T_3179_re;
    _T_3180_im <= _T_3179_im;
    _T_3181_re <= _T_3180_re;
    _T_3181_im <= _T_3180_im;
    _T_3182_re <= _T_3181_re;
    _T_3182_im <= _T_3181_im;
    _T_3183_re <= _T_3182_re;
    _T_3183_im <= _T_3182_im;
    _T_3184_re <= _T_3183_re;
    _T_3184_im <= _T_3183_im;
    _T_3185_re <= _T_3184_re;
    _T_3185_im <= _T_3184_im;
    _T_3186_re <= _T_3185_re;
    _T_3186_im <= _T_3185_im;
    _T_3187_re <= _T_3186_re;
    _T_3187_im <= _T_3186_im;
    _T_3188_re <= _T_3187_re;
    _T_3188_im <= _T_3187_im;
    _T_3189_re <= _T_3188_re;
    _T_3189_im <= _T_3188_im;
    _T_3190_re <= _T_3189_re;
    _T_3190_im <= _T_3189_im;
    _T_3191_re <= _T_3190_re;
    _T_3191_im <= _T_3190_im;
    _T_3192_re <= _T_3191_re;
    _T_3192_im <= _T_3191_im;
    _T_3193_re <= _T_3192_re;
    _T_3193_im <= _T_3192_im;
    _T_3194_re <= _T_3193_re;
    _T_3194_im <= _T_3193_im;
    _T_3195_re <= _T_3194_re;
    _T_3195_im <= _T_3194_im;
    _T_3196_re <= _T_3195_re;
    _T_3196_im <= _T_3195_im;
    _T_3197_re <= _T_3196_re;
    _T_3197_im <= _T_3196_im;
    _T_3198_re <= _T_3197_re;
    _T_3198_im <= _T_3197_im;
    _T_3199_re <= _T_3198_re;
    _T_3199_im <= _T_3198_im;
    _T_3200_re <= _T_3199_re;
    _T_3200_im <= _T_3199_im;
    _T_3201_re <= _T_3200_re;
    _T_3201_im <= _T_3200_im;
    _T_3202_re <= _T_3201_re;
    _T_3202_im <= _T_3201_im;
    _T_3203_re <= _T_3202_re;
    _T_3203_im <= _T_3202_im;
    _T_3204_re <= _T_3203_re;
    _T_3204_im <= _T_3203_im;
    _T_3205_re <= _T_3204_re;
    _T_3205_im <= _T_3204_im;
    _T_3206_re <= _T_3205_re;
    _T_3206_im <= _T_3205_im;
    _T_3207_re <= _T_3206_re;
    _T_3207_im <= _T_3206_im;
    _T_3208_re <= _T_3207_re;
    _T_3208_im <= _T_3207_im;
    _T_3209_re <= _T_3208_re;
    _T_3209_im <= _T_3208_im;
    _T_3210_re <= _T_3209_re;
    _T_3210_im <= _T_3209_im;
    _T_3211_re <= _T_3210_re;
    _T_3211_im <= _T_3210_im;
    _T_3212_re <= _T_3211_re;
    _T_3212_im <= _T_3211_im;
    _T_3213_re <= _T_3212_re;
    _T_3213_im <= _T_3212_im;
    _T_3214_re <= _T_3213_re;
    _T_3214_im <= _T_3213_im;
    _T_3215_re <= _T_3214_re;
    _T_3215_im <= _T_3214_im;
    _T_3216_re <= _T_3215_re;
    _T_3216_im <= _T_3215_im;
    _T_3217_re <= _T_3216_re;
    _T_3217_im <= _T_3216_im;
    _T_3218_re <= _T_3217_re;
    _T_3218_im <= _T_3217_im;
    _T_3219_re <= _T_3218_re;
    _T_3219_im <= _T_3218_im;
    _T_3220_re <= _T_3219_re;
    _T_3220_im <= _T_3219_im;
    _T_3221_re <= _T_3220_re;
    _T_3221_im <= _T_3220_im;
    _T_3222_re <= _T_3221_re;
    _T_3222_im <= _T_3221_im;
    _T_3223_re <= _T_3222_re;
    _T_3223_im <= _T_3222_im;
    _T_3224_re <= _T_3223_re;
    _T_3224_im <= _T_3223_im;
    _T_3225_re <= _T_3224_re;
    _T_3225_im <= _T_3224_im;
    _T_3226_re <= _T_3225_re;
    _T_3226_im <= _T_3225_im;
    _T_3227_re <= _T_3226_re;
    _T_3227_im <= _T_3226_im;
    _T_3228_re <= _T_3227_re;
    _T_3228_im <= _T_3227_im;
    _T_3229_re <= _T_3228_re;
    _T_3229_im <= _T_3228_im;
    _T_3230_re <= _T_3229_re;
    _T_3230_im <= _T_3229_im;
    _T_3231_re <= _T_3230_re;
    _T_3231_im <= _T_3230_im;
    _T_3232_re <= _T_3231_re;
    _T_3232_im <= _T_3231_im;
    _T_3233_re <= _T_3232_re;
    _T_3233_im <= _T_3232_im;
    _T_3234_re <= _T_3233_re;
    _T_3234_im <= _T_3233_im;
    _T_3235_re <= _T_3234_re;
    _T_3235_im <= _T_3234_im;
    _T_3236_re <= _T_3235_re;
    _T_3236_im <= _T_3235_im;
    _T_3237_re <= _T_3236_re;
    _T_3237_im <= _T_3236_im;
    _T_3238_re <= _T_3237_re;
    _T_3238_im <= _T_3237_im;
    _T_3239_re <= _T_3238_re;
    _T_3239_im <= _T_3238_im;
    _T_3240_re <= _T_3239_re;
    _T_3240_im <= _T_3239_im;
    _T_3241_re <= _T_3240_re;
    _T_3241_im <= _T_3240_im;
    _T_3242_re <= _T_3241_re;
    _T_3242_im <= _T_3241_im;
    _T_3243_re <= _T_3242_re;
    _T_3243_im <= _T_3242_im;
    _T_3244_re <= _T_3243_re;
    _T_3244_im <= _T_3243_im;
    _T_3245_re <= _T_3244_re;
    _T_3245_im <= _T_3244_im;
    _T_3246_re <= _T_3245_re;
    _T_3246_im <= _T_3245_im;
    _T_3247_re <= _T_3246_re;
    _T_3247_im <= _T_3246_im;
    _T_3248_re <= _T_3247_re;
    _T_3248_im <= _T_3247_im;
    _T_3249_re <= _T_3248_re;
    _T_3249_im <= _T_3248_im;
    _T_3250_re <= _T_3249_re;
    _T_3250_im <= _T_3249_im;
    _T_3251_re <= _T_3250_re;
    _T_3251_im <= _T_3250_im;
    _T_3252_re <= _T_3251_re;
    _T_3252_im <= _T_3251_im;
    _T_3253_re <= _T_3252_re;
    _T_3253_im <= _T_3252_im;
    _T_3254_re <= _T_3253_re;
    _T_3254_im <= _T_3253_im;
    _T_3255_re <= _T_3254_re;
    _T_3255_im <= _T_3254_im;
    _T_3256_re <= _T_3255_re;
    _T_3256_im <= _T_3255_im;
    _T_3257_re <= _T_3256_re;
    _T_3257_im <= _T_3256_im;
    _T_3258_re <= _T_3257_re;
    _T_3258_im <= _T_3257_im;
    _T_3259_re <= _T_3258_re;
    _T_3259_im <= _T_3258_im;
    _T_3260_re <= _T_3259_re;
    _T_3260_im <= _T_3259_im;
    _T_3261_re <= _T_3260_re;
    _T_3261_im <= _T_3260_im;
    _T_3262_re <= _T_3261_re;
    _T_3262_im <= _T_3261_im;
    _T_3268_re <= Switch_io_out1_re;
    _T_3268_im <= Switch_io_out1_im;
    _T_3269_re <= _T_3268_re;
    _T_3269_im <= _T_3268_im;
    _T_3270_re <= _T_3269_re;
    _T_3270_im <= _T_3269_im;
    _T_3271_re <= _T_3270_re;
    _T_3271_im <= _T_3270_im;
    _T_3272_re <= _T_3271_re;
    _T_3272_im <= _T_3271_im;
    _T_3273_re <= _T_3272_re;
    _T_3273_im <= _T_3272_im;
    _T_3274_re <= _T_3273_re;
    _T_3274_im <= _T_3273_im;
    _T_3275_re <= _T_3274_re;
    _T_3275_im <= _T_3274_im;
    _T_3276_re <= _T_3275_re;
    _T_3276_im <= _T_3275_im;
    _T_3277_re <= _T_3276_re;
    _T_3277_im <= _T_3276_im;
    _T_3278_re <= _T_3277_re;
    _T_3278_im <= _T_3277_im;
    _T_3279_re <= _T_3278_re;
    _T_3279_im <= _T_3278_im;
    _T_3280_re <= _T_3279_re;
    _T_3280_im <= _T_3279_im;
    _T_3281_re <= _T_3280_re;
    _T_3281_im <= _T_3280_im;
    _T_3282_re <= _T_3281_re;
    _T_3282_im <= _T_3281_im;
    _T_3283_re <= _T_3282_re;
    _T_3283_im <= _T_3282_im;
    _T_3284_re <= _T_3283_re;
    _T_3284_im <= _T_3283_im;
    _T_3285_re <= _T_3284_re;
    _T_3285_im <= _T_3284_im;
    _T_3286_re <= _T_3285_re;
    _T_3286_im <= _T_3285_im;
    _T_3287_re <= _T_3286_re;
    _T_3287_im <= _T_3286_im;
    _T_3288_re <= _T_3287_re;
    _T_3288_im <= _T_3287_im;
    _T_3289_re <= _T_3288_re;
    _T_3289_im <= _T_3288_im;
    _T_3290_re <= _T_3289_re;
    _T_3290_im <= _T_3289_im;
    _T_3291_re <= _T_3290_re;
    _T_3291_im <= _T_3290_im;
    _T_3292_re <= _T_3291_re;
    _T_3292_im <= _T_3291_im;
    _T_3293_re <= _T_3292_re;
    _T_3293_im <= _T_3292_im;
    _T_3294_re <= _T_3293_re;
    _T_3294_im <= _T_3293_im;
    _T_3295_re <= _T_3294_re;
    _T_3295_im <= _T_3294_im;
    _T_3296_re <= _T_3295_re;
    _T_3296_im <= _T_3295_im;
    _T_3297_re <= _T_3296_re;
    _T_3297_im <= _T_3296_im;
    _T_3298_re <= _T_3297_re;
    _T_3298_im <= _T_3297_im;
    _T_3299_re <= _T_3298_re;
    _T_3299_im <= _T_3298_im;
    _T_3300_re <= _T_3299_re;
    _T_3300_im <= _T_3299_im;
    _T_3301_re <= _T_3300_re;
    _T_3301_im <= _T_3300_im;
    _T_3302_re <= _T_3301_re;
    _T_3302_im <= _T_3301_im;
    _T_3303_re <= _T_3302_re;
    _T_3303_im <= _T_3302_im;
    _T_3304_re <= _T_3303_re;
    _T_3304_im <= _T_3303_im;
    _T_3305_re <= _T_3304_re;
    _T_3305_im <= _T_3304_im;
    _T_3306_re <= _T_3305_re;
    _T_3306_im <= _T_3305_im;
    _T_3307_re <= _T_3306_re;
    _T_3307_im <= _T_3306_im;
    _T_3308_re <= _T_3307_re;
    _T_3308_im <= _T_3307_im;
    _T_3309_re <= _T_3308_re;
    _T_3309_im <= _T_3308_im;
    _T_3310_re <= _T_3309_re;
    _T_3310_im <= _T_3309_im;
    _T_3311_re <= _T_3310_re;
    _T_3311_im <= _T_3310_im;
    _T_3312_re <= _T_3311_re;
    _T_3312_im <= _T_3311_im;
    _T_3313_re <= _T_3312_re;
    _T_3313_im <= _T_3312_im;
    _T_3314_re <= _T_3313_re;
    _T_3314_im <= _T_3313_im;
    _T_3315_re <= _T_3314_re;
    _T_3315_im <= _T_3314_im;
    _T_3316_re <= _T_3315_re;
    _T_3316_im <= _T_3315_im;
    _T_3317_re <= _T_3316_re;
    _T_3317_im <= _T_3316_im;
    _T_3318_re <= _T_3317_re;
    _T_3318_im <= _T_3317_im;
    _T_3319_re <= _T_3318_re;
    _T_3319_im <= _T_3318_im;
    _T_3320_re <= _T_3319_re;
    _T_3320_im <= _T_3319_im;
    _T_3321_re <= _T_3320_re;
    _T_3321_im <= _T_3320_im;
    _T_3322_re <= _T_3321_re;
    _T_3322_im <= _T_3321_im;
    _T_3323_re <= _T_3322_re;
    _T_3323_im <= _T_3322_im;
    _T_3324_re <= _T_3323_re;
    _T_3324_im <= _T_3323_im;
    _T_3325_re <= _T_3324_re;
    _T_3325_im <= _T_3324_im;
    _T_3326_re <= _T_3325_re;
    _T_3326_im <= _T_3325_im;
    _T_3327_re <= _T_3326_re;
    _T_3327_im <= _T_3326_im;
    _T_3328_re <= _T_3327_re;
    _T_3328_im <= _T_3327_im;
    _T_3329_re <= _T_3328_re;
    _T_3329_im <= _T_3328_im;
    _T_3330_re <= _T_3329_re;
    _T_3330_im <= _T_3329_im;
    _T_3331_re <= _T_3330_re;
    _T_3331_im <= _T_3330_im;
    _T_3332_re <= _T_3331_re;
    _T_3332_im <= _T_3331_im;
    _T_3333_re <= _T_3332_re;
    _T_3333_im <= _T_3332_im;
    _T_3334_re <= _T_3333_re;
    _T_3334_im <= _T_3333_im;
    _T_3335_re <= _T_3334_re;
    _T_3335_im <= _T_3334_im;
    _T_3336_re <= _T_3335_re;
    _T_3336_im <= _T_3335_im;
    _T_3337_re <= _T_3336_re;
    _T_3337_im <= _T_3336_im;
    _T_3338_re <= _T_3337_re;
    _T_3338_im <= _T_3337_im;
    _T_3339_re <= _T_3338_re;
    _T_3339_im <= _T_3338_im;
    _T_3340_re <= _T_3339_re;
    _T_3340_im <= _T_3339_im;
    _T_3341_re <= _T_3340_re;
    _T_3341_im <= _T_3340_im;
    _T_3342_re <= _T_3341_re;
    _T_3342_im <= _T_3341_im;
    _T_3343_re <= _T_3342_re;
    _T_3343_im <= _T_3342_im;
    _T_3344_re <= _T_3343_re;
    _T_3344_im <= _T_3343_im;
    _T_3345_re <= _T_3344_re;
    _T_3345_im <= _T_3344_im;
    _T_3346_re <= _T_3345_re;
    _T_3346_im <= _T_3345_im;
    _T_3347_re <= _T_3346_re;
    _T_3347_im <= _T_3346_im;
    _T_3348_re <= _T_3347_re;
    _T_3348_im <= _T_3347_im;
    _T_3349_re <= _T_3348_re;
    _T_3349_im <= _T_3348_im;
    _T_3350_re <= _T_3349_re;
    _T_3350_im <= _T_3349_im;
    _T_3351_re <= _T_3350_re;
    _T_3351_im <= _T_3350_im;
    _T_3352_re <= _T_3351_re;
    _T_3352_im <= _T_3351_im;
    _T_3353_re <= _T_3352_re;
    _T_3353_im <= _T_3352_im;
    _T_3354_re <= _T_3353_re;
    _T_3354_im <= _T_3353_im;
    _T_3355_re <= _T_3354_re;
    _T_3355_im <= _T_3354_im;
    _T_3356_re <= _T_3355_re;
    _T_3356_im <= _T_3355_im;
    _T_3357_re <= _T_3356_re;
    _T_3357_im <= _T_3356_im;
    _T_3358_re <= _T_3357_re;
    _T_3358_im <= _T_3357_im;
    _T_3359_re <= _T_3358_re;
    _T_3359_im <= _T_3358_im;
    _T_3360_re <= _T_3359_re;
    _T_3360_im <= _T_3359_im;
    _T_3361_re <= _T_3360_re;
    _T_3361_im <= _T_3360_im;
    _T_3362_re <= _T_3361_re;
    _T_3362_im <= _T_3361_im;
    _T_3363_re <= _T_3362_re;
    _T_3363_im <= _T_3362_im;
    _T_3364_re <= _T_3363_re;
    _T_3364_im <= _T_3363_im;
    _T_3365_re <= _T_3364_re;
    _T_3365_im <= _T_3364_im;
    _T_3366_re <= _T_3365_re;
    _T_3366_im <= _T_3365_im;
    _T_3367_re <= _T_3366_re;
    _T_3367_im <= _T_3366_im;
    _T_3368_re <= _T_3367_re;
    _T_3368_im <= _T_3367_im;
    _T_3369_re <= _T_3368_re;
    _T_3369_im <= _T_3368_im;
    _T_3370_re <= _T_3369_re;
    _T_3370_im <= _T_3369_im;
    _T_3371_re <= _T_3370_re;
    _T_3371_im <= _T_3370_im;
    _T_3372_re <= _T_3371_re;
    _T_3372_im <= _T_3371_im;
    _T_3373_re <= _T_3372_re;
    _T_3373_im <= _T_3372_im;
    _T_3374_re <= _T_3373_re;
    _T_3374_im <= _T_3373_im;
    _T_3375_re <= _T_3374_re;
    _T_3375_im <= _T_3374_im;
    _T_3376_re <= _T_3375_re;
    _T_3376_im <= _T_3375_im;
    _T_3377_re <= _T_3376_re;
    _T_3377_im <= _T_3376_im;
    _T_3378_re <= _T_3377_re;
    _T_3378_im <= _T_3377_im;
    _T_3379_re <= _T_3378_re;
    _T_3379_im <= _T_3378_im;
    _T_3380_re <= _T_3379_re;
    _T_3380_im <= _T_3379_im;
    _T_3381_re <= _T_3380_re;
    _T_3381_im <= _T_3380_im;
    _T_3382_re <= _T_3381_re;
    _T_3382_im <= _T_3381_im;
    _T_3383_re <= _T_3382_re;
    _T_3383_im <= _T_3382_im;
    _T_3384_re <= _T_3383_re;
    _T_3384_im <= _T_3383_im;
    _T_3385_re <= _T_3384_re;
    _T_3385_im <= _T_3384_im;
    _T_3386_re <= _T_3385_re;
    _T_3386_im <= _T_3385_im;
    _T_3387_re <= _T_3386_re;
    _T_3387_im <= _T_3386_im;
    _T_3388_re <= _T_3387_re;
    _T_3388_im <= _T_3387_im;
    _T_3389_re <= _T_3388_re;
    _T_3389_im <= _T_3388_im;
    _T_3390_re <= _T_3389_re;
    _T_3390_im <= _T_3389_im;
    _T_3391_re <= _T_3390_re;
    _T_3391_im <= _T_3390_im;
    _T_3392_re <= _T_3391_re;
    _T_3392_im <= _T_3391_im;
    _T_3393_re <= _T_3392_re;
    _T_3393_im <= _T_3392_im;
    _T_3394_re <= _T_3393_re;
    _T_3394_im <= _T_3393_im;
    _T_3395_re <= _T_3394_re;
    _T_3395_im <= _T_3394_im;
    _T_3396_re <= _T_3395_re;
    _T_3396_im <= _T_3395_im;
    _T_3397_re <= _T_3396_re;
    _T_3397_im <= _T_3396_im;
    _T_3398_re <= _T_3397_re;
    _T_3398_im <= _T_3397_im;
    _T_3399_re <= _T_3398_re;
    _T_3399_im <= _T_3398_im;
    _T_3400_re <= _T_3399_re;
    _T_3400_im <= _T_3399_im;
    _T_3401_re <= _T_3400_re;
    _T_3401_im <= _T_3400_im;
    _T_3402_re <= _T_3401_re;
    _T_3402_im <= _T_3401_im;
    _T_3403_re <= _T_3402_re;
    _T_3403_im <= _T_3402_im;
    _T_3404_re <= _T_3403_re;
    _T_3404_im <= _T_3403_im;
    _T_3405_re <= _T_3404_re;
    _T_3405_im <= _T_3404_im;
    _T_3406_re <= _T_3405_re;
    _T_3406_im <= _T_3405_im;
    _T_3407_re <= _T_3406_re;
    _T_3407_im <= _T_3406_im;
    _T_3408_re <= _T_3407_re;
    _T_3408_im <= _T_3407_im;
    _T_3409_re <= _T_3408_re;
    _T_3409_im <= _T_3408_im;
    _T_3410_re <= _T_3409_re;
    _T_3410_im <= _T_3409_im;
    _T_3411_re <= _T_3410_re;
    _T_3411_im <= _T_3410_im;
    _T_3412_re <= _T_3411_re;
    _T_3412_im <= _T_3411_im;
    _T_3413_re <= _T_3412_re;
    _T_3413_im <= _T_3412_im;
    _T_3414_re <= _T_3413_re;
    _T_3414_im <= _T_3413_im;
    _T_3415_re <= _T_3414_re;
    _T_3415_im <= _T_3414_im;
    _T_3416_re <= _T_3415_re;
    _T_3416_im <= _T_3415_im;
    _T_3417_re <= _T_3416_re;
    _T_3417_im <= _T_3416_im;
    _T_3418_re <= _T_3417_re;
    _T_3418_im <= _T_3417_im;
    _T_3419_re <= _T_3418_re;
    _T_3419_im <= _T_3418_im;
    _T_3420_re <= _T_3419_re;
    _T_3420_im <= _T_3419_im;
    _T_3421_re <= _T_3420_re;
    _T_3421_im <= _T_3420_im;
    _T_3422_re <= _T_3421_re;
    _T_3422_im <= _T_3421_im;
    _T_3423_re <= _T_3422_re;
    _T_3423_im <= _T_3422_im;
    _T_3424_re <= _T_3423_re;
    _T_3424_im <= _T_3423_im;
    _T_3425_re <= _T_3424_re;
    _T_3425_im <= _T_3424_im;
    _T_3426_re <= _T_3425_re;
    _T_3426_im <= _T_3425_im;
    _T_3427_re <= _T_3426_re;
    _T_3427_im <= _T_3426_im;
    _T_3428_re <= _T_3427_re;
    _T_3428_im <= _T_3427_im;
    _T_3429_re <= _T_3428_re;
    _T_3429_im <= _T_3428_im;
    _T_3430_re <= _T_3429_re;
    _T_3430_im <= _T_3429_im;
    _T_3431_re <= _T_3430_re;
    _T_3431_im <= _T_3430_im;
    _T_3432_re <= _T_3431_re;
    _T_3432_im <= _T_3431_im;
    _T_3433_re <= _T_3432_re;
    _T_3433_im <= _T_3432_im;
    _T_3434_re <= _T_3433_re;
    _T_3434_im <= _T_3433_im;
    _T_3435_re <= _T_3434_re;
    _T_3435_im <= _T_3434_im;
    _T_3436_re <= _T_3435_re;
    _T_3436_im <= _T_3435_im;
    _T_3437_re <= _T_3436_re;
    _T_3437_im <= _T_3436_im;
    _T_3438_re <= _T_3437_re;
    _T_3438_im <= _T_3437_im;
    _T_3439_re <= _T_3438_re;
    _T_3439_im <= _T_3438_im;
    _T_3440_re <= _T_3439_re;
    _T_3440_im <= _T_3439_im;
    _T_3441_re <= _T_3440_re;
    _T_3441_im <= _T_3440_im;
    _T_3442_re <= _T_3441_re;
    _T_3442_im <= _T_3441_im;
    _T_3443_re <= _T_3442_re;
    _T_3443_im <= _T_3442_im;
    _T_3444_re <= _T_3443_re;
    _T_3444_im <= _T_3443_im;
    _T_3445_re <= _T_3444_re;
    _T_3445_im <= _T_3444_im;
    _T_3446_re <= _T_3445_re;
    _T_3446_im <= _T_3445_im;
    _T_3447_re <= _T_3446_re;
    _T_3447_im <= _T_3446_im;
    _T_3448_re <= _T_3447_re;
    _T_3448_im <= _T_3447_im;
    _T_3449_re <= _T_3448_re;
    _T_3449_im <= _T_3448_im;
    _T_3450_re <= _T_3449_re;
    _T_3450_im <= _T_3449_im;
    _T_3451_re <= _T_3450_re;
    _T_3451_im <= _T_3450_im;
    _T_3452_re <= _T_3451_re;
    _T_3452_im <= _T_3451_im;
    _T_3453_re <= _T_3452_re;
    _T_3453_im <= _T_3452_im;
    _T_3454_re <= _T_3453_re;
    _T_3454_im <= _T_3453_im;
    _T_3455_re <= _T_3454_re;
    _T_3455_im <= _T_3454_im;
    _T_3456_re <= _T_3455_re;
    _T_3456_im <= _T_3455_im;
    _T_3457_re <= _T_3456_re;
    _T_3457_im <= _T_3456_im;
    _T_3458_re <= _T_3457_re;
    _T_3458_im <= _T_3457_im;
    _T_3459_re <= _T_3458_re;
    _T_3459_im <= _T_3458_im;
    _T_3460_re <= _T_3459_re;
    _T_3460_im <= _T_3459_im;
    _T_3461_re <= _T_3460_re;
    _T_3461_im <= _T_3460_im;
    _T_3462_re <= _T_3461_re;
    _T_3462_im <= _T_3461_im;
    _T_3463_re <= _T_3462_re;
    _T_3463_im <= _T_3462_im;
    _T_3464_re <= _T_3463_re;
    _T_3464_im <= _T_3463_im;
    _T_3465_re <= _T_3464_re;
    _T_3465_im <= _T_3464_im;
    _T_3466_re <= _T_3465_re;
    _T_3466_im <= _T_3465_im;
    _T_3467_re <= _T_3466_re;
    _T_3467_im <= _T_3466_im;
    _T_3468_re <= _T_3467_re;
    _T_3468_im <= _T_3467_im;
    _T_3469_re <= _T_3468_re;
    _T_3469_im <= _T_3468_im;
    _T_3470_re <= _T_3469_re;
    _T_3470_im <= _T_3469_im;
    _T_3471_re <= _T_3470_re;
    _T_3471_im <= _T_3470_im;
    _T_3472_re <= _T_3471_re;
    _T_3472_im <= _T_3471_im;
    _T_3473_re <= _T_3472_re;
    _T_3473_im <= _T_3472_im;
    _T_3474_re <= _T_3473_re;
    _T_3474_im <= _T_3473_im;
    _T_3475_re <= _T_3474_re;
    _T_3475_im <= _T_3474_im;
    _T_3476_re <= _T_3475_re;
    _T_3476_im <= _T_3475_im;
    _T_3477_re <= _T_3476_re;
    _T_3477_im <= _T_3476_im;
    _T_3478_re <= _T_3477_re;
    _T_3478_im <= _T_3477_im;
    _T_3479_re <= _T_3478_re;
    _T_3479_im <= _T_3478_im;
    _T_3480_re <= _T_3479_re;
    _T_3480_im <= _T_3479_im;
    _T_3481_re <= _T_3480_re;
    _T_3481_im <= _T_3480_im;
    _T_3482_re <= _T_3481_re;
    _T_3482_im <= _T_3481_im;
    _T_3483_re <= _T_3482_re;
    _T_3483_im <= _T_3482_im;
    _T_3484_re <= _T_3483_re;
    _T_3484_im <= _T_3483_im;
    _T_3485_re <= _T_3484_re;
    _T_3485_im <= _T_3484_im;
    _T_3486_re <= _T_3485_re;
    _T_3486_im <= _T_3485_im;
    _T_3487_re <= _T_3486_re;
    _T_3487_im <= _T_3486_im;
    _T_3488_re <= _T_3487_re;
    _T_3488_im <= _T_3487_im;
    _T_3489_re <= _T_3488_re;
    _T_3489_im <= _T_3488_im;
    _T_3490_re <= _T_3489_re;
    _T_3490_im <= _T_3489_im;
    _T_3491_re <= _T_3490_re;
    _T_3491_im <= _T_3490_im;
    _T_3492_re <= _T_3491_re;
    _T_3492_im <= _T_3491_im;
    _T_3493_re <= _T_3492_re;
    _T_3493_im <= _T_3492_im;
    _T_3494_re <= _T_3493_re;
    _T_3494_im <= _T_3493_im;
    _T_3495_re <= _T_3494_re;
    _T_3495_im <= _T_3494_im;
    _T_3496_re <= _T_3495_re;
    _T_3496_im <= _T_3495_im;
    _T_3497_re <= _T_3496_re;
    _T_3497_im <= _T_3496_im;
    _T_3498_re <= _T_3497_re;
    _T_3498_im <= _T_3497_im;
    _T_3499_re <= _T_3498_re;
    _T_3499_im <= _T_3498_im;
    _T_3500_re <= _T_3499_re;
    _T_3500_im <= _T_3499_im;
    _T_3501_re <= _T_3500_re;
    _T_3501_im <= _T_3500_im;
    _T_3502_re <= _T_3501_re;
    _T_3502_im <= _T_3501_im;
    _T_3503_re <= _T_3502_re;
    _T_3503_im <= _T_3502_im;
    _T_3504_re <= _T_3503_re;
    _T_3504_im <= _T_3503_im;
    _T_3505_re <= _T_3504_re;
    _T_3505_im <= _T_3504_im;
    _T_3506_re <= _T_3505_re;
    _T_3506_im <= _T_3505_im;
    _T_3507_re <= _T_3506_re;
    _T_3507_im <= _T_3506_im;
    _T_3508_re <= _T_3507_re;
    _T_3508_im <= _T_3507_im;
    _T_3509_re <= _T_3508_re;
    _T_3509_im <= _T_3508_im;
    _T_3510_re <= _T_3509_re;
    _T_3510_im <= _T_3509_im;
    _T_3511_re <= _T_3510_re;
    _T_3511_im <= _T_3510_im;
    _T_3512_re <= _T_3511_re;
    _T_3512_im <= _T_3511_im;
    _T_3513_re <= _T_3512_re;
    _T_3513_im <= _T_3512_im;
    _T_3514_re <= _T_3513_re;
    _T_3514_im <= _T_3513_im;
    _T_3515_re <= _T_3514_re;
    _T_3515_im <= _T_3514_im;
    _T_3516_re <= _T_3515_re;
    _T_3516_im <= _T_3515_im;
    _T_3517_re <= _T_3516_re;
    _T_3517_im <= _T_3516_im;
    _T_3518_re <= _T_3517_re;
    _T_3518_im <= _T_3517_im;
    _T_3519_re <= _T_3518_re;
    _T_3519_im <= _T_3518_im;
    _T_3520_re <= _T_3519_re;
    _T_3520_im <= _T_3519_im;
    _T_3521_re <= _T_3520_re;
    _T_3521_im <= _T_3520_im;
    _T_3522_re <= _T_3521_re;
    _T_3522_im <= _T_3521_im;
    _T_3523_re <= _T_3522_re;
    _T_3523_im <= _T_3522_im;
    _T_3524_re <= _T_3523_re;
    _T_3524_im <= _T_3523_im;
    _T_3525_re <= _T_3524_re;
    _T_3525_im <= _T_3524_im;
    _T_3526_re <= _T_3525_re;
    _T_3526_im <= _T_3525_im;
    _T_3527_re <= _T_3526_re;
    _T_3527_im <= _T_3526_im;
    _T_3528_re <= _T_3527_re;
    _T_3528_im <= _T_3527_im;
    _T_3529_re <= _T_3528_re;
    _T_3529_im <= _T_3528_im;
    _T_3530_re <= _T_3529_re;
    _T_3530_im <= _T_3529_im;
    _T_3531_re <= _T_3530_re;
    _T_3531_im <= _T_3530_im;
    _T_3532_re <= _T_3531_re;
    _T_3532_im <= _T_3531_im;
    _T_3533_re <= _T_3532_re;
    _T_3533_im <= _T_3532_im;
    _T_3534_re <= _T_3533_re;
    _T_3534_im <= _T_3533_im;
    _T_3535_re <= _T_3534_re;
    _T_3535_im <= _T_3534_im;
    _T_3536_re <= _T_3535_re;
    _T_3536_im <= _T_3535_im;
    _T_3537_re <= _T_3536_re;
    _T_3537_im <= _T_3536_im;
    _T_3538_re <= _T_3537_re;
    _T_3538_im <= _T_3537_im;
    _T_3539_re <= _T_3538_re;
    _T_3539_im <= _T_3538_im;
    _T_3540_re <= _T_3539_re;
    _T_3540_im <= _T_3539_im;
    _T_3541_re <= _T_3540_re;
    _T_3541_im <= _T_3540_im;
    _T_3542_re <= _T_3541_re;
    _T_3542_im <= _T_3541_im;
    _T_3543_re <= _T_3542_re;
    _T_3543_im <= _T_3542_im;
    _T_3544_re <= _T_3543_re;
    _T_3544_im <= _T_3543_im;
    _T_3545_re <= _T_3544_re;
    _T_3545_im <= _T_3544_im;
    _T_3546_re <= _T_3545_re;
    _T_3546_im <= _T_3545_im;
    _T_3547_re <= _T_3546_re;
    _T_3547_im <= _T_3546_im;
    _T_3548_re <= _T_3547_re;
    _T_3548_im <= _T_3547_im;
    _T_3549_re <= _T_3548_re;
    _T_3549_im <= _T_3548_im;
    _T_3550_re <= _T_3549_re;
    _T_3550_im <= _T_3549_im;
    _T_3551_re <= _T_3550_re;
    _T_3551_im <= _T_3550_im;
    _T_3552_re <= _T_3551_re;
    _T_3552_im <= _T_3551_im;
    _T_3553_re <= _T_3552_re;
    _T_3553_im <= _T_3552_im;
    _T_3554_re <= _T_3553_re;
    _T_3554_im <= _T_3553_im;
    _T_3555_re <= _T_3554_re;
    _T_3555_im <= _T_3554_im;
    _T_3556_re <= _T_3555_re;
    _T_3556_im <= _T_3555_im;
    _T_3557_re <= _T_3556_re;
    _T_3557_im <= _T_3556_im;
    _T_3558_re <= _T_3557_re;
    _T_3558_im <= _T_3557_im;
    _T_3559_re <= _T_3558_re;
    _T_3559_im <= _T_3558_im;
    _T_3560_re <= _T_3559_re;
    _T_3560_im <= _T_3559_im;
    _T_3561_re <= _T_3560_re;
    _T_3561_im <= _T_3560_im;
    _T_3562_re <= _T_3561_re;
    _T_3562_im <= _T_3561_im;
    _T_3563_re <= _T_3562_re;
    _T_3563_im <= _T_3562_im;
    _T_3564_re <= _T_3563_re;
    _T_3564_im <= _T_3563_im;
    _T_3565_re <= _T_3564_re;
    _T_3565_im <= _T_3564_im;
    _T_3566_re <= _T_3565_re;
    _T_3566_im <= _T_3565_im;
    _T_3567_re <= _T_3566_re;
    _T_3567_im <= _T_3566_im;
    _T_3568_re <= _T_3567_re;
    _T_3568_im <= _T_3567_im;
    _T_3569_re <= _T_3568_re;
    _T_3569_im <= _T_3568_im;
    _T_3570_re <= _T_3569_re;
    _T_3570_im <= _T_3569_im;
    _T_3571_re <= _T_3570_re;
    _T_3571_im <= _T_3570_im;
    _T_3572_re <= _T_3571_re;
    _T_3572_im <= _T_3571_im;
    _T_3573_re <= _T_3572_re;
    _T_3573_im <= _T_3572_im;
    _T_3574_re <= _T_3573_re;
    _T_3574_im <= _T_3573_im;
    _T_3575_re <= _T_3574_re;
    _T_3575_im <= _T_3574_im;
    _T_3576_re <= _T_3575_re;
    _T_3576_im <= _T_3575_im;
    _T_3577_re <= _T_3576_re;
    _T_3577_im <= _T_3576_im;
    _T_3578_re <= _T_3577_re;
    _T_3578_im <= _T_3577_im;
    _T_3579_re <= _T_3578_re;
    _T_3579_im <= _T_3578_im;
    _T_3580_re <= _T_3579_re;
    _T_3580_im <= _T_3579_im;
    _T_3581_re <= _T_3580_re;
    _T_3581_im <= _T_3580_im;
    _T_3582_re <= _T_3581_re;
    _T_3582_im <= _T_3581_im;
    _T_3583_re <= _T_3582_re;
    _T_3583_im <= _T_3582_im;
    _T_3584_re <= _T_3583_re;
    _T_3584_im <= _T_3583_im;
    _T_3585_re <= _T_3584_re;
    _T_3585_im <= _T_3584_im;
    _T_3586_re <= _T_3585_re;
    _T_3586_im <= _T_3585_im;
    _T_3587_re <= _T_3586_re;
    _T_3587_im <= _T_3586_im;
    _T_3588_re <= _T_3587_re;
    _T_3588_im <= _T_3587_im;
    _T_3589_re <= _T_3588_re;
    _T_3589_im <= _T_3588_im;
    _T_3590_re <= _T_3589_re;
    _T_3590_im <= _T_3589_im;
    _T_3591_re <= _T_3590_re;
    _T_3591_im <= _T_3590_im;
    _T_3592_re <= _T_3591_re;
    _T_3592_im <= _T_3591_im;
    _T_3593_re <= _T_3592_re;
    _T_3593_im <= _T_3592_im;
    _T_3594_re <= _T_3593_re;
    _T_3594_im <= _T_3593_im;
    _T_3595_re <= _T_3594_re;
    _T_3595_im <= _T_3594_im;
    _T_3596_re <= _T_3595_re;
    _T_3596_im <= _T_3595_im;
    _T_3597_re <= _T_3596_re;
    _T_3597_im <= _T_3596_im;
    _T_3598_re <= _T_3597_re;
    _T_3598_im <= _T_3597_im;
    _T_3599_re <= _T_3598_re;
    _T_3599_im <= _T_3598_im;
    _T_3600_re <= _T_3599_re;
    _T_3600_im <= _T_3599_im;
    _T_3601_re <= _T_3600_re;
    _T_3601_im <= _T_3600_im;
    _T_3602_re <= _T_3601_re;
    _T_3602_im <= _T_3601_im;
    _T_3603_re <= _T_3602_re;
    _T_3603_im <= _T_3602_im;
    _T_3604_re <= _T_3603_re;
    _T_3604_im <= _T_3603_im;
    _T_3605_re <= _T_3604_re;
    _T_3605_im <= _T_3604_im;
    _T_3606_re <= _T_3605_re;
    _T_3606_im <= _T_3605_im;
    _T_3607_re <= _T_3606_re;
    _T_3607_im <= _T_3606_im;
    _T_3608_re <= _T_3607_re;
    _T_3608_im <= _T_3607_im;
    _T_3609_re <= _T_3608_re;
    _T_3609_im <= _T_3608_im;
    _T_3610_re <= _T_3609_re;
    _T_3610_im <= _T_3609_im;
    _T_3611_re <= _T_3610_re;
    _T_3611_im <= _T_3610_im;
    _T_3612_re <= _T_3611_re;
    _T_3612_im <= _T_3611_im;
    _T_3613_re <= _T_3612_re;
    _T_3613_im <= _T_3612_im;
    _T_3614_re <= _T_3613_re;
    _T_3614_im <= _T_3613_im;
    _T_3615_re <= _T_3614_re;
    _T_3615_im <= _T_3614_im;
    _T_3616_re <= _T_3615_re;
    _T_3616_im <= _T_3615_im;
    _T_3617_re <= _T_3616_re;
    _T_3617_im <= _T_3616_im;
    _T_3618_re <= _T_3617_re;
    _T_3618_im <= _T_3617_im;
    _T_3619_re <= _T_3618_re;
    _T_3619_im <= _T_3618_im;
    _T_3620_re <= _T_3619_re;
    _T_3620_im <= _T_3619_im;
    _T_3621_re <= _T_3620_re;
    _T_3621_im <= _T_3620_im;
    _T_3622_re <= _T_3621_re;
    _T_3622_im <= _T_3621_im;
    _T_3623_re <= _T_3622_re;
    _T_3623_im <= _T_3622_im;
    _T_3624_re <= _T_3623_re;
    _T_3624_im <= _T_3623_im;
    _T_3625_re <= _T_3624_re;
    _T_3625_im <= _T_3624_im;
    _T_3626_re <= _T_3625_re;
    _T_3626_im <= _T_3625_im;
    _T_3627_re <= _T_3626_re;
    _T_3627_im <= _T_3626_im;
    _T_3628_re <= _T_3627_re;
    _T_3628_im <= _T_3627_im;
    _T_3629_re <= _T_3628_re;
    _T_3629_im <= _T_3628_im;
    _T_3630_re <= _T_3629_re;
    _T_3630_im <= _T_3629_im;
    _T_3631_re <= _T_3630_re;
    _T_3631_im <= _T_3630_im;
    _T_3632_re <= _T_3631_re;
    _T_3632_im <= _T_3631_im;
    _T_3633_re <= _T_3632_re;
    _T_3633_im <= _T_3632_im;
    _T_3634_re <= _T_3633_re;
    _T_3634_im <= _T_3633_im;
    _T_3635_re <= _T_3634_re;
    _T_3635_im <= _T_3634_im;
    _T_3636_re <= _T_3635_re;
    _T_3636_im <= _T_3635_im;
    _T_3637_re <= _T_3636_re;
    _T_3637_im <= _T_3636_im;
    _T_3638_re <= _T_3637_re;
    _T_3638_im <= _T_3637_im;
    _T_3639_re <= _T_3638_re;
    _T_3639_im <= _T_3638_im;
    _T_3640_re <= _T_3639_re;
    _T_3640_im <= _T_3639_im;
    _T_3641_re <= _T_3640_re;
    _T_3641_im <= _T_3640_im;
    _T_3642_re <= _T_3641_re;
    _T_3642_im <= _T_3641_im;
    _T_3643_re <= _T_3642_re;
    _T_3643_im <= _T_3642_im;
    _T_3644_re <= _T_3643_re;
    _T_3644_im <= _T_3643_im;
    _T_3645_re <= _T_3644_re;
    _T_3645_im <= _T_3644_im;
    _T_3646_re <= _T_3645_re;
    _T_3646_im <= _T_3645_im;
    _T_3647_re <= _T_3646_re;
    _T_3647_im <= _T_3646_im;
    _T_3648_re <= _T_3647_re;
    _T_3648_im <= _T_3647_im;
    _T_3649_re <= _T_3648_re;
    _T_3649_im <= _T_3648_im;
    _T_3650_re <= _T_3649_re;
    _T_3650_im <= _T_3649_im;
    _T_3651_re <= _T_3650_re;
    _T_3651_im <= _T_3650_im;
    _T_3652_re <= _T_3651_re;
    _T_3652_im <= _T_3651_im;
    _T_3653_re <= _T_3652_re;
    _T_3653_im <= _T_3652_im;
    _T_3654_re <= _T_3653_re;
    _T_3654_im <= _T_3653_im;
    _T_3655_re <= _T_3654_re;
    _T_3655_im <= _T_3654_im;
    _T_3656_re <= _T_3655_re;
    _T_3656_im <= _T_3655_im;
    _T_3657_re <= _T_3656_re;
    _T_3657_im <= _T_3656_im;
    _T_3658_re <= _T_3657_re;
    _T_3658_im <= _T_3657_im;
    _T_3659_re <= _T_3658_re;
    _T_3659_im <= _T_3658_im;
    _T_3660_re <= _T_3659_re;
    _T_3660_im <= _T_3659_im;
    _T_3661_re <= _T_3660_re;
    _T_3661_im <= _T_3660_im;
    _T_3662_re <= _T_3661_re;
    _T_3662_im <= _T_3661_im;
    _T_3663_re <= _T_3662_re;
    _T_3663_im <= _T_3662_im;
    _T_3664_re <= _T_3663_re;
    _T_3664_im <= _T_3663_im;
    _T_3665_re <= _T_3664_re;
    _T_3665_im <= _T_3664_im;
    _T_3666_re <= _T_3665_re;
    _T_3666_im <= _T_3665_im;
    _T_3667_re <= _T_3666_re;
    _T_3667_im <= _T_3666_im;
    _T_3668_re <= _T_3667_re;
    _T_3668_im <= _T_3667_im;
    _T_3669_re <= _T_3668_re;
    _T_3669_im <= _T_3668_im;
    _T_3670_re <= _T_3669_re;
    _T_3670_im <= _T_3669_im;
    _T_3671_re <= _T_3670_re;
    _T_3671_im <= _T_3670_im;
    _T_3672_re <= _T_3671_re;
    _T_3672_im <= _T_3671_im;
    _T_3673_re <= _T_3672_re;
    _T_3673_im <= _T_3672_im;
    _T_3674_re <= _T_3673_re;
    _T_3674_im <= _T_3673_im;
    _T_3675_re <= _T_3674_re;
    _T_3675_im <= _T_3674_im;
    _T_3676_re <= _T_3675_re;
    _T_3676_im <= _T_3675_im;
    _T_3677_re <= _T_3676_re;
    _T_3677_im <= _T_3676_im;
    _T_3678_re <= _T_3677_re;
    _T_3678_im <= _T_3677_im;
    _T_3679_re <= _T_3678_re;
    _T_3679_im <= _T_3678_im;
    _T_3680_re <= _T_3679_re;
    _T_3680_im <= _T_3679_im;
    _T_3681_re <= _T_3680_re;
    _T_3681_im <= _T_3680_im;
    _T_3682_re <= _T_3681_re;
    _T_3682_im <= _T_3681_im;
    _T_3683_re <= _T_3682_re;
    _T_3683_im <= _T_3682_im;
    _T_3684_re <= _T_3683_re;
    _T_3684_im <= _T_3683_im;
    _T_3685_re <= _T_3684_re;
    _T_3685_im <= _T_3684_im;
    _T_3686_re <= _T_3685_re;
    _T_3686_im <= _T_3685_im;
    _T_3687_re <= _T_3686_re;
    _T_3687_im <= _T_3686_im;
    _T_3688_re <= _T_3687_re;
    _T_3688_im <= _T_3687_im;
    _T_3689_re <= _T_3688_re;
    _T_3689_im <= _T_3688_im;
    _T_3690_re <= _T_3689_re;
    _T_3690_im <= _T_3689_im;
    _T_3691_re <= _T_3690_re;
    _T_3691_im <= _T_3690_im;
    _T_3692_re <= _T_3691_re;
    _T_3692_im <= _T_3691_im;
    _T_3693_re <= _T_3692_re;
    _T_3693_im <= _T_3692_im;
    _T_3694_re <= _T_3693_re;
    _T_3694_im <= _T_3693_im;
    _T_3695_re <= _T_3694_re;
    _T_3695_im <= _T_3694_im;
    _T_3696_re <= _T_3695_re;
    _T_3696_im <= _T_3695_im;
    _T_3697_re <= _T_3696_re;
    _T_3697_im <= _T_3696_im;
    _T_3698_re <= _T_3697_re;
    _T_3698_im <= _T_3697_im;
    _T_3699_re <= _T_3698_re;
    _T_3699_im <= _T_3698_im;
    _T_3700_re <= _T_3699_re;
    _T_3700_im <= _T_3699_im;
    _T_3701_re <= _T_3700_re;
    _T_3701_im <= _T_3700_im;
    _T_3702_re <= _T_3701_re;
    _T_3702_im <= _T_3701_im;
    _T_3703_re <= _T_3702_re;
    _T_3703_im <= _T_3702_im;
    _T_3704_re <= _T_3703_re;
    _T_3704_im <= _T_3703_im;
    _T_3705_re <= _T_3704_re;
    _T_3705_im <= _T_3704_im;
    _T_3706_re <= _T_3705_re;
    _T_3706_im <= _T_3705_im;
    _T_3707_re <= _T_3706_re;
    _T_3707_im <= _T_3706_im;
    _T_3708_re <= _T_3707_re;
    _T_3708_im <= _T_3707_im;
    _T_3709_re <= _T_3708_re;
    _T_3709_im <= _T_3708_im;
    _T_3710_re <= _T_3709_re;
    _T_3710_im <= _T_3709_im;
    _T_3711_re <= _T_3710_re;
    _T_3711_im <= _T_3710_im;
    _T_3712_re <= _T_3711_re;
    _T_3712_im <= _T_3711_im;
    _T_3713_re <= _T_3712_re;
    _T_3713_im <= _T_3712_im;
    _T_3714_re <= _T_3713_re;
    _T_3714_im <= _T_3713_im;
    _T_3715_re <= _T_3714_re;
    _T_3715_im <= _T_3714_im;
    _T_3716_re <= _T_3715_re;
    _T_3716_im <= _T_3715_im;
    _T_3717_re <= _T_3716_re;
    _T_3717_im <= _T_3716_im;
    _T_3718_re <= _T_3717_re;
    _T_3718_im <= _T_3717_im;
    _T_3719_re <= _T_3718_re;
    _T_3719_im <= _T_3718_im;
    _T_3720_re <= _T_3719_re;
    _T_3720_im <= _T_3719_im;
    _T_3721_re <= _T_3720_re;
    _T_3721_im <= _T_3720_im;
    _T_3722_re <= _T_3721_re;
    _T_3722_im <= _T_3721_im;
    _T_3723_re <= _T_3722_re;
    _T_3723_im <= _T_3722_im;
    _T_3724_re <= _T_3723_re;
    _T_3724_im <= _T_3723_im;
    _T_3725_re <= _T_3724_re;
    _T_3725_im <= _T_3724_im;
    _T_3726_re <= _T_3725_re;
    _T_3726_im <= _T_3725_im;
    _T_3727_re <= _T_3726_re;
    _T_3727_im <= _T_3726_im;
    _T_3728_re <= _T_3727_re;
    _T_3728_im <= _T_3727_im;
    _T_3729_re <= _T_3728_re;
    _T_3729_im <= _T_3728_im;
    _T_3730_re <= _T_3729_re;
    _T_3730_im <= _T_3729_im;
    _T_3731_re <= _T_3730_re;
    _T_3731_im <= _T_3730_im;
    _T_3732_re <= _T_3731_re;
    _T_3732_im <= _T_3731_im;
    _T_3733_re <= _T_3732_re;
    _T_3733_im <= _T_3732_im;
    _T_3734_re <= _T_3733_re;
    _T_3734_im <= _T_3733_im;
    _T_3735_re <= _T_3734_re;
    _T_3735_im <= _T_3734_im;
    _T_3736_re <= _T_3735_re;
    _T_3736_im <= _T_3735_im;
    _T_3737_re <= _T_3736_re;
    _T_3737_im <= _T_3736_im;
    _T_3738_re <= _T_3737_re;
    _T_3738_im <= _T_3737_im;
    _T_3739_re <= _T_3738_re;
    _T_3739_im <= _T_3738_im;
    _T_3740_re <= _T_3739_re;
    _T_3740_im <= _T_3739_im;
    _T_3741_re <= _T_3740_re;
    _T_3741_im <= _T_3740_im;
    _T_3742_re <= _T_3741_re;
    _T_3742_im <= _T_3741_im;
    _T_3743_re <= _T_3742_re;
    _T_3743_im <= _T_3742_im;
    _T_3744_re <= _T_3743_re;
    _T_3744_im <= _T_3743_im;
    _T_3745_re <= _T_3744_re;
    _T_3745_im <= _T_3744_im;
    _T_3746_re <= _T_3745_re;
    _T_3746_im <= _T_3745_im;
    _T_3747_re <= _T_3746_re;
    _T_3747_im <= _T_3746_im;
    _T_3748_re <= _T_3747_re;
    _T_3748_im <= _T_3747_im;
    _T_3749_re <= _T_3748_re;
    _T_3749_im <= _T_3748_im;
    _T_3750_re <= _T_3749_re;
    _T_3750_im <= _T_3749_im;
    _T_3751_re <= _T_3750_re;
    _T_3751_im <= _T_3750_im;
    _T_3752_re <= _T_3751_re;
    _T_3752_im <= _T_3751_im;
    _T_3753_re <= _T_3752_re;
    _T_3753_im <= _T_3752_im;
    _T_3754_re <= _T_3753_re;
    _T_3754_im <= _T_3753_im;
    _T_3755_re <= _T_3754_re;
    _T_3755_im <= _T_3754_im;
    _T_3756_re <= _T_3755_re;
    _T_3756_im <= _T_3755_im;
    _T_3757_re <= _T_3756_re;
    _T_3757_im <= _T_3756_im;
    _T_3758_re <= _T_3757_re;
    _T_3758_im <= _T_3757_im;
    _T_3759_re <= _T_3758_re;
    _T_3759_im <= _T_3758_im;
    _T_3760_re <= _T_3759_re;
    _T_3760_im <= _T_3759_im;
    _T_3761_re <= _T_3760_re;
    _T_3761_im <= _T_3760_im;
    _T_3762_re <= _T_3761_re;
    _T_3762_im <= _T_3761_im;
    _T_3763_re <= _T_3762_re;
    _T_3763_im <= _T_3762_im;
    _T_3764_re <= _T_3763_re;
    _T_3764_im <= _T_3763_im;
    _T_3765_re <= _T_3764_re;
    _T_3765_im <= _T_3764_im;
    _T_3766_re <= _T_3765_re;
    _T_3766_im <= _T_3765_im;
    _T_3767_re <= _T_3766_re;
    _T_3767_im <= _T_3766_im;
    _T_3768_re <= _T_3767_re;
    _T_3768_im <= _T_3767_im;
    _T_3769_re <= _T_3768_re;
    _T_3769_im <= _T_3768_im;
    _T_3770_re <= _T_3769_re;
    _T_3770_im <= _T_3769_im;
    _T_3771_re <= _T_3770_re;
    _T_3771_im <= _T_3770_im;
    _T_3772_re <= _T_3771_re;
    _T_3772_im <= _T_3771_im;
    _T_3773_re <= _T_3772_re;
    _T_3773_im <= _T_3772_im;
    _T_3774_re <= _T_3773_re;
    _T_3774_im <= _T_3773_im;
    _T_3775_re <= _T_3774_re;
    _T_3775_im <= _T_3774_im;
    _T_3776_re <= _T_3775_re;
    _T_3776_im <= _T_3775_im;
    _T_3777_re <= _T_3776_re;
    _T_3777_im <= _T_3776_im;
    _T_3778_re <= _T_3777_re;
    _T_3778_im <= _T_3777_im;
    _T_3779_re <= _T_3778_re;
    _T_3779_im <= _T_3778_im;
    _T_3780_re <= _T_3779_re;
    _T_3780_im <= _T_3779_im;
    _T_3781_re <= _T_3780_re;
    _T_3781_im <= _T_3780_im;
    _T_3782_re <= _T_3781_re;
    _T_3782_im <= _T_3781_im;
    _T_3783_re <= _T_3782_re;
    _T_3783_im <= _T_3782_im;
    _T_3784_re <= _T_3783_re;
    _T_3784_im <= _T_3783_im;
    _T_3785_re <= _T_3784_re;
    _T_3785_im <= _T_3784_im;
    _T_3786_re <= _T_3785_re;
    _T_3786_im <= _T_3785_im;
    _T_3787_re <= _T_3786_re;
    _T_3787_im <= _T_3786_im;
    _T_3788_re <= _T_3787_re;
    _T_3788_im <= _T_3787_im;
    _T_3789_re <= _T_3788_re;
    _T_3789_im <= _T_3788_im;
    _T_3790_re <= _T_3789_re;
    _T_3790_im <= _T_3789_im;
    _T_3791_re <= _T_3790_re;
    _T_3791_im <= _T_3790_im;
    _T_3792_re <= _T_3791_re;
    _T_3792_im <= _T_3791_im;
    _T_3793_re <= _T_3792_re;
    _T_3793_im <= _T_3792_im;
    _T_3794_re <= _T_3793_re;
    _T_3794_im <= _T_3793_im;
    _T_3795_re <= _T_3794_re;
    _T_3795_im <= _T_3794_im;
    _T_3796_re <= _T_3795_re;
    _T_3796_im <= _T_3795_im;
    _T_3797_re <= _T_3796_re;
    _T_3797_im <= _T_3796_im;
    _T_3798_re <= _T_3797_re;
    _T_3798_im <= _T_3797_im;
    _T_3799_re <= _T_3798_re;
    _T_3799_im <= _T_3798_im;
    _T_3800_re <= _T_3799_re;
    _T_3800_im <= _T_3799_im;
    _T_3801_re <= _T_3800_re;
    _T_3801_im <= _T_3800_im;
    _T_3802_re <= _T_3801_re;
    _T_3802_im <= _T_3801_im;
    _T_3803_re <= _T_3802_re;
    _T_3803_im <= _T_3802_im;
    _T_3804_re <= _T_3803_re;
    _T_3804_im <= _T_3803_im;
    _T_3805_re <= _T_3804_re;
    _T_3805_im <= _T_3804_im;
    _T_3806_re <= _T_3805_re;
    _T_3806_im <= _T_3805_im;
    _T_3807_re <= _T_3806_re;
    _T_3807_im <= _T_3806_im;
    _T_3808_re <= _T_3807_re;
    _T_3808_im <= _T_3807_im;
    _T_3809_re <= _T_3808_re;
    _T_3809_im <= _T_3808_im;
    _T_3810_re <= _T_3809_re;
    _T_3810_im <= _T_3809_im;
    _T_3811_re <= _T_3810_re;
    _T_3811_im <= _T_3810_im;
    _T_3812_re <= _T_3811_re;
    _T_3812_im <= _T_3811_im;
    _T_3813_re <= _T_3812_re;
    _T_3813_im <= _T_3812_im;
    _T_3814_re <= _T_3813_re;
    _T_3814_im <= _T_3813_im;
    _T_3815_re <= _T_3814_re;
    _T_3815_im <= _T_3814_im;
    _T_3816_re <= _T_3815_re;
    _T_3816_im <= _T_3815_im;
    _T_3817_re <= _T_3816_re;
    _T_3817_im <= _T_3816_im;
    _T_3818_re <= _T_3817_re;
    _T_3818_im <= _T_3817_im;
    _T_3819_re <= _T_3818_re;
    _T_3819_im <= _T_3818_im;
    _T_3820_re <= _T_3819_re;
    _T_3820_im <= _T_3819_im;
    _T_3821_re <= _T_3820_re;
    _T_3821_im <= _T_3820_im;
    _T_3822_re <= _T_3821_re;
    _T_3822_im <= _T_3821_im;
    _T_3823_re <= _T_3822_re;
    _T_3823_im <= _T_3822_im;
    _T_3824_re <= _T_3823_re;
    _T_3824_im <= _T_3823_im;
    _T_3825_re <= _T_3824_re;
    _T_3825_im <= _T_3824_im;
    _T_3826_re <= _T_3825_re;
    _T_3826_im <= _T_3825_im;
    _T_3827_re <= _T_3826_re;
    _T_3827_im <= _T_3826_im;
    _T_3828_re <= _T_3827_re;
    _T_3828_im <= _T_3827_im;
    _T_3829_re <= _T_3828_re;
    _T_3829_im <= _T_3828_im;
    _T_3830_re <= _T_3829_re;
    _T_3830_im <= _T_3829_im;
    _T_3831_re <= _T_3830_re;
    _T_3831_im <= _T_3830_im;
    _T_3832_re <= _T_3831_re;
    _T_3832_im <= _T_3831_im;
    _T_3833_re <= _T_3832_re;
    _T_3833_im <= _T_3832_im;
    _T_3834_re <= _T_3833_re;
    _T_3834_im <= _T_3833_im;
    _T_3835_re <= _T_3834_re;
    _T_3835_im <= _T_3834_im;
    _T_3836_re <= _T_3835_re;
    _T_3836_im <= _T_3835_im;
    _T_3837_re <= _T_3836_re;
    _T_3837_im <= _T_3836_im;
    _T_3838_re <= _T_3837_re;
    _T_3838_im <= _T_3837_im;
    _T_3839_re <= _T_3838_re;
    _T_3839_im <= _T_3838_im;
    _T_3840_re <= _T_3839_re;
    _T_3840_im <= _T_3839_im;
    _T_3841_re <= _T_3840_re;
    _T_3841_im <= _T_3840_im;
    _T_3842_re <= _T_3841_re;
    _T_3842_im <= _T_3841_im;
    _T_3843_re <= _T_3842_re;
    _T_3843_im <= _T_3842_im;
    _T_3844_re <= _T_3843_re;
    _T_3844_im <= _T_3843_im;
    _T_3845_re <= _T_3844_re;
    _T_3845_im <= _T_3844_im;
    _T_3846_re <= _T_3845_re;
    _T_3846_im <= _T_3845_im;
    _T_3847_re <= _T_3846_re;
    _T_3847_im <= _T_3846_im;
    _T_3848_re <= _T_3847_re;
    _T_3848_im <= _T_3847_im;
    _T_3849_re <= _T_3848_re;
    _T_3849_im <= _T_3848_im;
    _T_3850_re <= _T_3849_re;
    _T_3850_im <= _T_3849_im;
    _T_3851_re <= _T_3850_re;
    _T_3851_im <= _T_3850_im;
    _T_3852_re <= _T_3851_re;
    _T_3852_im <= _T_3851_im;
    _T_3853_re <= _T_3852_re;
    _T_3853_im <= _T_3852_im;
    _T_3854_re <= _T_3853_re;
    _T_3854_im <= _T_3853_im;
    _T_3855_re <= _T_3854_re;
    _T_3855_im <= _T_3854_im;
    _T_3856_re <= _T_3855_re;
    _T_3856_im <= _T_3855_im;
    _T_3857_re <= _T_3856_re;
    _T_3857_im <= _T_3856_im;
    _T_3858_re <= _T_3857_re;
    _T_3858_im <= _T_3857_im;
    _T_3859_re <= _T_3858_re;
    _T_3859_im <= _T_3858_im;
    _T_3860_re <= _T_3859_re;
    _T_3860_im <= _T_3859_im;
    _T_3861_re <= _T_3860_re;
    _T_3861_im <= _T_3860_im;
    _T_3862_re <= _T_3861_re;
    _T_3862_im <= _T_3861_im;
    _T_3863_re <= _T_3862_re;
    _T_3863_im <= _T_3862_im;
    _T_3864_re <= _T_3863_re;
    _T_3864_im <= _T_3863_im;
    _T_3865_re <= _T_3864_re;
    _T_3865_im <= _T_3864_im;
    _T_3866_re <= _T_3865_re;
    _T_3866_im <= _T_3865_im;
    _T_3867_re <= _T_3866_re;
    _T_3867_im <= _T_3866_im;
    _T_3868_re <= _T_3867_re;
    _T_3868_im <= _T_3867_im;
    _T_3869_re <= _T_3868_re;
    _T_3869_im <= _T_3868_im;
    _T_3870_re <= _T_3869_re;
    _T_3870_im <= _T_3869_im;
    _T_3871_re <= _T_3870_re;
    _T_3871_im <= _T_3870_im;
    _T_3872_re <= _T_3871_re;
    _T_3872_im <= _T_3871_im;
    _T_3873_re <= _T_3872_re;
    _T_3873_im <= _T_3872_im;
    _T_3874_re <= _T_3873_re;
    _T_3874_im <= _T_3873_im;
    _T_3875_re <= _T_3874_re;
    _T_3875_im <= _T_3874_im;
    _T_3876_re <= _T_3875_re;
    _T_3876_im <= _T_3875_im;
    _T_3877_re <= _T_3876_re;
    _T_3877_im <= _T_3876_im;
    _T_3878_re <= _T_3877_re;
    _T_3878_im <= _T_3877_im;
    _T_3879_re <= _T_3878_re;
    _T_3879_im <= _T_3878_im;
    _T_3880_re <= _T_3879_re;
    _T_3880_im <= _T_3879_im;
    _T_3881_re <= _T_3880_re;
    _T_3881_im <= _T_3880_im;
    _T_3882_re <= _T_3881_re;
    _T_3882_im <= _T_3881_im;
    _T_3883_re <= _T_3882_re;
    _T_3883_im <= _T_3882_im;
    _T_3884_re <= _T_3883_re;
    _T_3884_im <= _T_3883_im;
    _T_3885_re <= _T_3884_re;
    _T_3885_im <= _T_3884_im;
    _T_3886_re <= _T_3885_re;
    _T_3886_im <= _T_3885_im;
    _T_3887_re <= _T_3886_re;
    _T_3887_im <= _T_3886_im;
    _T_3888_re <= _T_3887_re;
    _T_3888_im <= _T_3887_im;
    _T_3889_re <= _T_3888_re;
    _T_3889_im <= _T_3888_im;
    _T_3890_re <= _T_3889_re;
    _T_3890_im <= _T_3889_im;
    _T_3891_re <= _T_3890_re;
    _T_3891_im <= _T_3890_im;
    _T_3892_re <= _T_3891_re;
    _T_3892_im <= _T_3891_im;
    _T_3893_re <= _T_3892_re;
    _T_3893_im <= _T_3892_im;
    _T_3894_re <= _T_3893_re;
    _T_3894_im <= _T_3893_im;
    _T_3895_re <= _T_3894_re;
    _T_3895_im <= _T_3894_im;
    _T_3896_re <= _T_3895_re;
    _T_3896_im <= _T_3895_im;
    _T_3897_re <= _T_3896_re;
    _T_3897_im <= _T_3896_im;
    _T_3898_re <= _T_3897_re;
    _T_3898_im <= _T_3897_im;
    _T_3899_re <= _T_3898_re;
    _T_3899_im <= _T_3898_im;
    _T_3900_re <= _T_3899_re;
    _T_3900_im <= _T_3899_im;
    _T_3901_re <= _T_3900_re;
    _T_3901_im <= _T_3900_im;
    _T_3902_re <= _T_3901_re;
    _T_3902_im <= _T_3901_im;
    _T_3903_re <= _T_3902_re;
    _T_3903_im <= _T_3902_im;
    _T_3904_re <= _T_3903_re;
    _T_3904_im <= _T_3903_im;
    _T_3905_re <= _T_3904_re;
    _T_3905_im <= _T_3904_im;
    _T_3906_re <= _T_3905_re;
    _T_3906_im <= _T_3905_im;
    _T_3907_re <= _T_3906_re;
    _T_3907_im <= _T_3906_im;
    _T_3908_re <= _T_3907_re;
    _T_3908_im <= _T_3907_im;
    _T_3909_re <= _T_3908_re;
    _T_3909_im <= _T_3908_im;
    _T_3910_re <= _T_3909_re;
    _T_3910_im <= _T_3909_im;
    _T_3911_re <= _T_3910_re;
    _T_3911_im <= _T_3910_im;
    _T_3912_re <= _T_3911_re;
    _T_3912_im <= _T_3911_im;
    _T_3913_re <= _T_3912_re;
    _T_3913_im <= _T_3912_im;
    _T_3914_re <= _T_3913_re;
    _T_3914_im <= _T_3913_im;
    _T_3915_re <= _T_3914_re;
    _T_3915_im <= _T_3914_im;
    _T_3916_re <= _T_3915_re;
    _T_3916_im <= _T_3915_im;
    _T_3917_re <= _T_3916_re;
    _T_3917_im <= _T_3916_im;
    _T_3918_re <= _T_3917_re;
    _T_3918_im <= _T_3917_im;
    _T_3919_re <= _T_3918_re;
    _T_3919_im <= _T_3918_im;
    _T_3920_re <= _T_3919_re;
    _T_3920_im <= _T_3919_im;
    _T_3921_re <= _T_3920_re;
    _T_3921_im <= _T_3920_im;
    _T_3922_re <= _T_3921_re;
    _T_3922_im <= _T_3921_im;
    _T_3923_re <= _T_3922_re;
    _T_3923_im <= _T_3922_im;
    _T_3924_re <= _T_3923_re;
    _T_3924_im <= _T_3923_im;
    _T_3925_re <= _T_3924_re;
    _T_3925_im <= _T_3924_im;
    _T_3926_re <= _T_3925_re;
    _T_3926_im <= _T_3925_im;
    _T_3927_re <= _T_3926_re;
    _T_3927_im <= _T_3926_im;
    _T_3928_re <= _T_3927_re;
    _T_3928_im <= _T_3927_im;
    _T_3929_re <= _T_3928_re;
    _T_3929_im <= _T_3928_im;
    _T_3930_re <= _T_3929_re;
    _T_3930_im <= _T_3929_im;
    _T_3931_re <= _T_3930_re;
    _T_3931_im <= _T_3930_im;
    _T_3932_re <= _T_3931_re;
    _T_3932_im <= _T_3931_im;
    _T_3933_re <= _T_3932_re;
    _T_3933_im <= _T_3932_im;
    _T_3934_re <= _T_3933_re;
    _T_3934_im <= _T_3933_im;
    _T_3935_re <= _T_3934_re;
    _T_3935_im <= _T_3934_im;
    _T_3936_re <= _T_3935_re;
    _T_3936_im <= _T_3935_im;
    _T_3937_re <= _T_3936_re;
    _T_3937_im <= _T_3936_im;
    _T_3938_re <= _T_3937_re;
    _T_3938_im <= _T_3937_im;
    _T_3939_re <= _T_3938_re;
    _T_3939_im <= _T_3938_im;
    _T_3940_re <= _T_3939_re;
    _T_3940_im <= _T_3939_im;
    _T_3941_re <= _T_3940_re;
    _T_3941_im <= _T_3940_im;
    _T_3942_re <= _T_3941_re;
    _T_3942_im <= _T_3941_im;
    _T_3943_re <= _T_3942_re;
    _T_3943_im <= _T_3942_im;
    _T_3944_re <= _T_3943_re;
    _T_3944_im <= _T_3943_im;
    _T_3945_re <= _T_3944_re;
    _T_3945_im <= _T_3944_im;
    _T_3946_re <= _T_3945_re;
    _T_3946_im <= _T_3945_im;
    _T_3947_re <= _T_3946_re;
    _T_3947_im <= _T_3946_im;
    _T_3948_re <= _T_3947_re;
    _T_3948_im <= _T_3947_im;
    _T_3949_re <= _T_3948_re;
    _T_3949_im <= _T_3948_im;
    _T_3950_re <= _T_3949_re;
    _T_3950_im <= _T_3949_im;
    _T_3951_re <= _T_3950_re;
    _T_3951_im <= _T_3950_im;
    _T_3952_re <= _T_3951_re;
    _T_3952_im <= _T_3951_im;
    _T_3953_re <= _T_3952_re;
    _T_3953_im <= _T_3952_im;
    _T_3954_re <= _T_3953_re;
    _T_3954_im <= _T_3953_im;
    _T_3955_re <= _T_3954_re;
    _T_3955_im <= _T_3954_im;
    _T_3956_re <= _T_3955_re;
    _T_3956_im <= _T_3955_im;
    _T_3957_re <= _T_3956_re;
    _T_3957_im <= _T_3956_im;
    _T_3958_re <= _T_3957_re;
    _T_3958_im <= _T_3957_im;
    _T_3959_re <= _T_3958_re;
    _T_3959_im <= _T_3958_im;
    _T_3960_re <= _T_3959_re;
    _T_3960_im <= _T_3959_im;
    _T_3961_re <= _T_3960_re;
    _T_3961_im <= _T_3960_im;
    _T_3962_re <= _T_3961_re;
    _T_3962_im <= _T_3961_im;
    _T_3963_re <= _T_3962_re;
    _T_3963_im <= _T_3962_im;
    _T_3964_re <= _T_3963_re;
    _T_3964_im <= _T_3963_im;
    _T_3965_re <= _T_3964_re;
    _T_3965_im <= _T_3964_im;
    _T_3966_re <= _T_3965_re;
    _T_3966_im <= _T_3965_im;
    _T_3967_re <= _T_3966_re;
    _T_3967_im <= _T_3966_im;
    _T_3968_re <= _T_3967_re;
    _T_3968_im <= _T_3967_im;
    _T_3969_re <= _T_3968_re;
    _T_3969_im <= _T_3968_im;
    _T_3970_re <= _T_3969_re;
    _T_3970_im <= _T_3969_im;
    _T_3971_re <= _T_3970_re;
    _T_3971_im <= _T_3970_im;
    _T_3972_re <= _T_3971_re;
    _T_3972_im <= _T_3971_im;
    _T_3973_re <= _T_3972_re;
    _T_3973_im <= _T_3972_im;
    _T_3974_re <= _T_3973_re;
    _T_3974_im <= _T_3973_im;
    _T_3975_re <= _T_3974_re;
    _T_3975_im <= _T_3974_im;
    _T_3976_re <= _T_3975_re;
    _T_3976_im <= _T_3975_im;
    _T_3977_re <= _T_3976_re;
    _T_3977_im <= _T_3976_im;
    _T_3978_re <= _T_3977_re;
    _T_3978_im <= _T_3977_im;
    _T_3979_re <= _T_3978_re;
    _T_3979_im <= _T_3978_im;
    _T_3980_re <= _T_3979_re;
    _T_3980_im <= _T_3979_im;
    _T_3981_re <= _T_3980_re;
    _T_3981_im <= _T_3980_im;
    _T_3982_re <= _T_3981_re;
    _T_3982_im <= _T_3981_im;
    _T_3983_re <= _T_3982_re;
    _T_3983_im <= _T_3982_im;
    _T_3984_re <= _T_3983_re;
    _T_3984_im <= _T_3983_im;
    _T_3985_re <= _T_3984_re;
    _T_3985_im <= _T_3984_im;
    _T_3986_re <= _T_3985_re;
    _T_3986_im <= _T_3985_im;
    _T_3987_re <= _T_3986_re;
    _T_3987_im <= _T_3986_im;
    _T_3988_re <= _T_3987_re;
    _T_3988_im <= _T_3987_im;
    _T_3989_re <= _T_3988_re;
    _T_3989_im <= _T_3988_im;
    _T_3990_re <= _T_3989_re;
    _T_3990_im <= _T_3989_im;
    _T_3991_re <= _T_3990_re;
    _T_3991_im <= _T_3990_im;
    _T_3992_re <= _T_3991_re;
    _T_3992_im <= _T_3991_im;
    _T_3993_re <= _T_3992_re;
    _T_3993_im <= _T_3992_im;
    _T_3994_re <= _T_3993_re;
    _T_3994_im <= _T_3993_im;
    _T_3995_re <= _T_3994_re;
    _T_3995_im <= _T_3994_im;
    _T_3996_re <= _T_3995_re;
    _T_3996_im <= _T_3995_im;
    _T_3997_re <= _T_3996_re;
    _T_3997_im <= _T_3996_im;
    _T_3998_re <= _T_3997_re;
    _T_3998_im <= _T_3997_im;
    _T_3999_re <= _T_3998_re;
    _T_3999_im <= _T_3998_im;
    _T_4000_re <= _T_3999_re;
    _T_4000_im <= _T_3999_im;
    _T_4001_re <= _T_4000_re;
    _T_4001_im <= _T_4000_im;
    _T_4002_re <= _T_4001_re;
    _T_4002_im <= _T_4001_im;
    _T_4003_re <= _T_4002_re;
    _T_4003_im <= _T_4002_im;
    _T_4004_re <= _T_4003_re;
    _T_4004_im <= _T_4003_im;
    _T_4005_re <= _T_4004_re;
    _T_4005_im <= _T_4004_im;
    _T_4006_re <= _T_4005_re;
    _T_4006_im <= _T_4005_im;
    _T_4007_re <= _T_4006_re;
    _T_4007_im <= _T_4006_im;
    _T_4008_re <= _T_4007_re;
    _T_4008_im <= _T_4007_im;
    _T_4009_re <= _T_4008_re;
    _T_4009_im <= _T_4008_im;
    _T_4010_re <= _T_4009_re;
    _T_4010_im <= _T_4009_im;
    _T_4011_re <= _T_4010_re;
    _T_4011_im <= _T_4010_im;
    _T_4012_re <= _T_4011_re;
    _T_4012_im <= _T_4011_im;
    _T_4013_re <= _T_4012_re;
    _T_4013_im <= _T_4012_im;
    _T_4014_re <= _T_4013_re;
    _T_4014_im <= _T_4013_im;
    _T_4015_re <= _T_4014_re;
    _T_4015_im <= _T_4014_im;
    _T_4016_re <= _T_4015_re;
    _T_4016_im <= _T_4015_im;
    _T_4017_re <= _T_4016_re;
    _T_4017_im <= _T_4016_im;
    _T_4018_re <= _T_4017_re;
    _T_4018_im <= _T_4017_im;
    _T_4019_re <= _T_4018_re;
    _T_4019_im <= _T_4018_im;
    _T_4020_re <= _T_4019_re;
    _T_4020_im <= _T_4019_im;
    _T_4021_re <= _T_4020_re;
    _T_4021_im <= _T_4020_im;
    _T_4022_re <= _T_4021_re;
    _T_4022_im <= _T_4021_im;
    _T_4023_re <= _T_4022_re;
    _T_4023_im <= _T_4022_im;
    _T_4024_re <= _T_4023_re;
    _T_4024_im <= _T_4023_im;
    _T_4025_re <= _T_4024_re;
    _T_4025_im <= _T_4024_im;
    _T_4026_re <= _T_4025_re;
    _T_4026_im <= _T_4025_im;
    _T_4027_re <= _T_4026_re;
    _T_4027_im <= _T_4026_im;
    _T_4028_re <= _T_4027_re;
    _T_4028_im <= _T_4027_im;
    _T_4029_re <= _T_4028_re;
    _T_4029_im <= _T_4028_im;
    _T_4030_re <= _T_4029_re;
    _T_4030_im <= _T_4029_im;
    _T_4031_re <= _T_4030_re;
    _T_4031_im <= _T_4030_im;
    _T_4032_re <= _T_4031_re;
    _T_4032_im <= _T_4031_im;
    _T_4033_re <= _T_4032_re;
    _T_4033_im <= _T_4032_im;
    _T_4034_re <= _T_4033_re;
    _T_4034_im <= _T_4033_im;
    _T_4035_re <= _T_4034_re;
    _T_4035_im <= _T_4034_im;
    _T_4036_re <= _T_4035_re;
    _T_4036_im <= _T_4035_im;
    _T_4037_re <= _T_4036_re;
    _T_4037_im <= _T_4036_im;
    _T_4038_re <= _T_4037_re;
    _T_4038_im <= _T_4037_im;
    _T_4039_re <= _T_4038_re;
    _T_4039_im <= _T_4038_im;
    _T_4040_re <= _T_4039_re;
    _T_4040_im <= _T_4039_im;
    _T_4041_re <= _T_4040_re;
    _T_4041_im <= _T_4040_im;
    _T_4042_re <= _T_4041_re;
    _T_4042_im <= _T_4041_im;
    _T_4043_re <= _T_4042_re;
    _T_4043_im <= _T_4042_im;
    _T_4044_re <= _T_4043_re;
    _T_4044_im <= _T_4043_im;
    _T_4045_re <= _T_4044_re;
    _T_4045_im <= _T_4044_im;
    _T_4046_re <= _T_4045_re;
    _T_4046_im <= _T_4045_im;
    _T_4047_re <= _T_4046_re;
    _T_4047_im <= _T_4046_im;
    _T_4048_re <= _T_4047_re;
    _T_4048_im <= _T_4047_im;
    _T_4049_re <= _T_4048_re;
    _T_4049_im <= _T_4048_im;
    _T_4050_re <= _T_4049_re;
    _T_4050_im <= _T_4049_im;
    _T_4051_re <= _T_4050_re;
    _T_4051_im <= _T_4050_im;
    _T_4052_re <= _T_4051_re;
    _T_4052_im <= _T_4051_im;
    _T_4053_re <= _T_4052_re;
    _T_4053_im <= _T_4052_im;
    _T_4054_re <= _T_4053_re;
    _T_4054_im <= _T_4053_im;
    _T_4055_re <= _T_4054_re;
    _T_4055_im <= _T_4054_im;
    _T_4056_re <= _T_4055_re;
    _T_4056_im <= _T_4055_im;
    _T_4057_re <= _T_4056_re;
    _T_4057_im <= _T_4056_im;
    _T_4058_re <= _T_4057_re;
    _T_4058_im <= _T_4057_im;
    _T_4059_re <= _T_4058_re;
    _T_4059_im <= _T_4058_im;
    _T_4060_re <= _T_4059_re;
    _T_4060_im <= _T_4059_im;
    _T_4061_re <= _T_4060_re;
    _T_4061_im <= _T_4060_im;
    _T_4062_re <= _T_4061_re;
    _T_4062_im <= _T_4061_im;
    _T_4063_re <= _T_4062_re;
    _T_4063_im <= _T_4062_im;
    _T_4064_re <= _T_4063_re;
    _T_4064_im <= _T_4063_im;
    _T_4065_re <= _T_4064_re;
    _T_4065_im <= _T_4064_im;
    _T_4066_re <= _T_4065_re;
    _T_4066_im <= _T_4065_im;
    _T_4067_re <= _T_4066_re;
    _T_4067_im <= _T_4066_im;
    _T_4068_re <= _T_4067_re;
    _T_4068_im <= _T_4067_im;
    _T_4069_re <= _T_4068_re;
    _T_4069_im <= _T_4068_im;
    _T_4070_re <= _T_4069_re;
    _T_4070_im <= _T_4069_im;
    _T_4071_re <= _T_4070_re;
    _T_4071_im <= _T_4070_im;
    _T_4072_re <= _T_4071_re;
    _T_4072_im <= _T_4071_im;
    _T_4073_re <= _T_4072_re;
    _T_4073_im <= _T_4072_im;
    _T_4074_re <= _T_4073_re;
    _T_4074_im <= _T_4073_im;
    _T_4075_re <= _T_4074_re;
    _T_4075_im <= _T_4074_im;
    _T_4076_re <= _T_4075_re;
    _T_4076_im <= _T_4075_im;
    _T_4077_re <= _T_4076_re;
    _T_4077_im <= _T_4076_im;
    _T_4078_re <= _T_4077_re;
    _T_4078_im <= _T_4077_im;
    _T_4079_re <= _T_4078_re;
    _T_4079_im <= _T_4078_im;
    _T_4080_re <= _T_4079_re;
    _T_4080_im <= _T_4079_im;
    _T_4081_re <= _T_4080_re;
    _T_4081_im <= _T_4080_im;
    _T_4082_re <= _T_4081_re;
    _T_4082_im <= _T_4081_im;
    _T_4083_re <= _T_4082_re;
    _T_4083_im <= _T_4082_im;
    _T_4084_re <= _T_4083_re;
    _T_4084_im <= _T_4083_im;
    _T_4085_re <= _T_4084_re;
    _T_4085_im <= _T_4084_im;
    _T_4086_re <= _T_4085_re;
    _T_4086_im <= _T_4085_im;
    _T_4087_re <= _T_4086_re;
    _T_4087_im <= _T_4086_im;
    _T_4088_re <= _T_4087_re;
    _T_4088_im <= _T_4087_im;
    _T_4089_re <= _T_4088_re;
    _T_4089_im <= _T_4088_im;
    _T_4090_re <= _T_4089_re;
    _T_4090_im <= _T_4089_im;
    _T_4091_re <= _T_4090_re;
    _T_4091_im <= _T_4090_im;
    _T_4092_re <= _T_4091_re;
    _T_4092_im <= _T_4091_im;
    _T_4093_re <= _T_4092_re;
    _T_4093_im <= _T_4092_im;
    _T_4094_re <= _T_4093_re;
    _T_4094_im <= _T_4093_im;
    _T_4095_re <= _T_4094_re;
    _T_4095_im <= _T_4094_im;
    _T_4096_re <= _T_4095_re;
    _T_4096_im <= _T_4095_im;
    _T_4097_re <= _T_4096_re;
    _T_4097_im <= _T_4096_im;
    _T_4098_re <= _T_4097_re;
    _T_4098_im <= _T_4097_im;
    _T_4099_re <= _T_4098_re;
    _T_4099_im <= _T_4098_im;
    _T_4100_re <= _T_4099_re;
    _T_4100_im <= _T_4099_im;
    _T_4101_re <= _T_4100_re;
    _T_4101_im <= _T_4100_im;
    _T_4102_re <= _T_4101_re;
    _T_4102_im <= _T_4101_im;
    _T_4103_re <= _T_4102_re;
    _T_4103_im <= _T_4102_im;
    _T_4104_re <= _T_4103_re;
    _T_4104_im <= _T_4103_im;
    _T_4105_re <= _T_4104_re;
    _T_4105_im <= _T_4104_im;
    _T_4106_re <= _T_4105_re;
    _T_4106_im <= _T_4105_im;
    _T_4107_re <= _T_4106_re;
    _T_4107_im <= _T_4106_im;
    _T_4108_re <= _T_4107_re;
    _T_4108_im <= _T_4107_im;
    _T_4109_re <= _T_4108_re;
    _T_4109_im <= _T_4108_im;
    _T_4110_re <= _T_4109_re;
    _T_4110_im <= _T_4109_im;
    _T_4111_re <= _T_4110_re;
    _T_4111_im <= _T_4110_im;
    _T_4112_re <= _T_4111_re;
    _T_4112_im <= _T_4111_im;
    _T_4113_re <= _T_4112_re;
    _T_4113_im <= _T_4112_im;
    _T_4114_re <= _T_4113_re;
    _T_4114_im <= _T_4113_im;
    _T_4115_re <= _T_4114_re;
    _T_4115_im <= _T_4114_im;
    _T_4116_re <= _T_4115_re;
    _T_4116_im <= _T_4115_im;
    _T_4117_re <= _T_4116_re;
    _T_4117_im <= _T_4116_im;
    _T_4118_re <= _T_4117_re;
    _T_4118_im <= _T_4117_im;
    _T_4119_re <= _T_4118_re;
    _T_4119_im <= _T_4118_im;
    _T_4120_re <= _T_4119_re;
    _T_4120_im <= _T_4119_im;
    _T_4121_re <= _T_4120_re;
    _T_4121_im <= _T_4120_im;
    _T_4122_re <= _T_4121_re;
    _T_4122_im <= _T_4121_im;
    _T_4123_re <= _T_4122_re;
    _T_4123_im <= _T_4122_im;
    _T_4124_re <= _T_4123_re;
    _T_4124_im <= _T_4123_im;
    _T_4125_re <= _T_4124_re;
    _T_4125_im <= _T_4124_im;
    _T_4126_re <= _T_4125_re;
    _T_4126_im <= _T_4125_im;
    _T_4127_re <= _T_4126_re;
    _T_4127_im <= _T_4126_im;
    _T_4128_re <= _T_4127_re;
    _T_4128_im <= _T_4127_im;
    _T_4129_re <= _T_4128_re;
    _T_4129_im <= _T_4128_im;
    _T_4130_re <= _T_4129_re;
    _T_4130_im <= _T_4129_im;
    _T_4131_re <= _T_4130_re;
    _T_4131_im <= _T_4130_im;
    _T_4132_re <= _T_4131_re;
    _T_4132_im <= _T_4131_im;
    _T_4133_re <= _T_4132_re;
    _T_4133_im <= _T_4132_im;
    _T_4134_re <= _T_4133_re;
    _T_4134_im <= _T_4133_im;
    _T_4135_re <= _T_4134_re;
    _T_4135_im <= _T_4134_im;
    _T_4136_re <= _T_4135_re;
    _T_4136_im <= _T_4135_im;
    _T_4137_re <= _T_4136_re;
    _T_4137_im <= _T_4136_im;
    _T_4138_re <= _T_4137_re;
    _T_4138_im <= _T_4137_im;
    _T_4139_re <= _T_4138_re;
    _T_4139_im <= _T_4138_im;
    _T_4140_re <= _T_4139_re;
    _T_4140_im <= _T_4139_im;
    _T_4141_re <= _T_4140_re;
    _T_4141_im <= _T_4140_im;
    _T_4142_re <= _T_4141_re;
    _T_4142_im <= _T_4141_im;
    _T_4143_re <= _T_4142_re;
    _T_4143_im <= _T_4142_im;
    _T_4144_re <= _T_4143_re;
    _T_4144_im <= _T_4143_im;
    _T_4145_re <= _T_4144_re;
    _T_4145_im <= _T_4144_im;
    _T_4146_re <= _T_4145_re;
    _T_4146_im <= _T_4145_im;
    _T_4147_re <= _T_4146_re;
    _T_4147_im <= _T_4146_im;
    _T_4148_re <= _T_4147_re;
    _T_4148_im <= _T_4147_im;
    _T_4149_re <= _T_4148_re;
    _T_4149_im <= _T_4148_im;
    _T_4150_re <= _T_4149_re;
    _T_4150_im <= _T_4149_im;
    _T_4151_re <= _T_4150_re;
    _T_4151_im <= _T_4150_im;
    _T_4152_re <= _T_4151_re;
    _T_4152_im <= _T_4151_im;
    _T_4153_re <= _T_4152_re;
    _T_4153_im <= _T_4152_im;
    _T_4154_re <= _T_4153_re;
    _T_4154_im <= _T_4153_im;
    _T_4155_re <= _T_4154_re;
    _T_4155_im <= _T_4154_im;
    _T_4156_re <= _T_4155_re;
    _T_4156_im <= _T_4155_im;
    _T_4157_re <= _T_4156_re;
    _T_4157_im <= _T_4156_im;
    _T_4158_re <= _T_4157_re;
    _T_4158_im <= _T_4157_im;
    _T_4159_re <= _T_4158_re;
    _T_4159_im <= _T_4158_im;
    _T_4160_re <= _T_4159_re;
    _T_4160_im <= _T_4159_im;
    _T_4161_re <= _T_4160_re;
    _T_4161_im <= _T_4160_im;
    _T_4162_re <= _T_4161_re;
    _T_4162_im <= _T_4161_im;
    _T_4163_re <= _T_4162_re;
    _T_4163_im <= _T_4162_im;
    _T_4164_re <= _T_4163_re;
    _T_4164_im <= _T_4163_im;
    _T_4165_re <= _T_4164_re;
    _T_4165_im <= _T_4164_im;
    _T_4166_re <= _T_4165_re;
    _T_4166_im <= _T_4165_im;
    _T_4167_re <= _T_4166_re;
    _T_4167_im <= _T_4166_im;
    _T_4168_re <= _T_4167_re;
    _T_4168_im <= _T_4167_im;
    _T_4169_re <= _T_4168_re;
    _T_4169_im <= _T_4168_im;
    _T_4170_re <= _T_4169_re;
    _T_4170_im <= _T_4169_im;
    _T_4171_re <= _T_4170_re;
    _T_4171_im <= _T_4170_im;
    _T_4172_re <= _T_4171_re;
    _T_4172_im <= _T_4171_im;
    _T_4173_re <= _T_4172_re;
    _T_4173_im <= _T_4172_im;
    _T_4174_re <= _T_4173_re;
    _T_4174_im <= _T_4173_im;
    _T_4175_re <= _T_4174_re;
    _T_4175_im <= _T_4174_im;
    _T_4176_re <= _T_4175_re;
    _T_4176_im <= _T_4175_im;
    _T_4177_re <= _T_4176_re;
    _T_4177_im <= _T_4176_im;
    _T_4178_re <= _T_4177_re;
    _T_4178_im <= _T_4177_im;
    _T_4179_re <= _T_4178_re;
    _T_4179_im <= _T_4178_im;
    _T_4180_re <= _T_4179_re;
    _T_4180_im <= _T_4179_im;
    _T_4181_re <= _T_4180_re;
    _T_4181_im <= _T_4180_im;
    _T_4182_re <= _T_4181_re;
    _T_4182_im <= _T_4181_im;
    _T_4183_re <= _T_4182_re;
    _T_4183_im <= _T_4182_im;
    _T_4184_re <= _T_4183_re;
    _T_4184_im <= _T_4183_im;
    _T_4185_re <= _T_4184_re;
    _T_4185_im <= _T_4184_im;
    _T_4186_re <= _T_4185_re;
    _T_4186_im <= _T_4185_im;
    _T_4187_re <= _T_4186_re;
    _T_4187_im <= _T_4186_im;
    _T_4188_re <= _T_4187_re;
    _T_4188_im <= _T_4187_im;
    _T_4189_re <= _T_4188_re;
    _T_4189_im <= _T_4188_im;
    _T_4190_re <= _T_4189_re;
    _T_4190_im <= _T_4189_im;
    _T_4191_re <= _T_4190_re;
    _T_4191_im <= _T_4190_im;
    _T_4192_re <= _T_4191_re;
    _T_4192_im <= _T_4191_im;
    _T_4193_re <= _T_4192_re;
    _T_4193_im <= _T_4192_im;
    _T_4194_re <= _T_4193_re;
    _T_4194_im <= _T_4193_im;
    _T_4195_re <= _T_4194_re;
    _T_4195_im <= _T_4194_im;
    _T_4196_re <= _T_4195_re;
    _T_4196_im <= _T_4195_im;
    _T_4197_re <= _T_4196_re;
    _T_4197_im <= _T_4196_im;
    _T_4198_re <= _T_4197_re;
    _T_4198_im <= _T_4197_im;
    _T_4199_re <= _T_4198_re;
    _T_4199_im <= _T_4198_im;
    _T_4200_re <= _T_4199_re;
    _T_4200_im <= _T_4199_im;
    _T_4201_re <= _T_4200_re;
    _T_4201_im <= _T_4200_im;
    _T_4202_re <= _T_4201_re;
    _T_4202_im <= _T_4201_im;
    _T_4203_re <= _T_4202_re;
    _T_4203_im <= _T_4202_im;
    _T_4204_re <= _T_4203_re;
    _T_4204_im <= _T_4203_im;
    _T_4205_re <= _T_4204_re;
    _T_4205_im <= _T_4204_im;
    _T_4206_re <= _T_4205_re;
    _T_4206_im <= _T_4205_im;
    _T_4207_re <= _T_4206_re;
    _T_4207_im <= _T_4206_im;
    _T_4208_re <= _T_4207_re;
    _T_4208_im <= _T_4207_im;
    _T_4209_re <= _T_4208_re;
    _T_4209_im <= _T_4208_im;
    _T_4210_re <= _T_4209_re;
    _T_4210_im <= _T_4209_im;
    _T_4211_re <= _T_4210_re;
    _T_4211_im <= _T_4210_im;
    _T_4212_re <= _T_4211_re;
    _T_4212_im <= _T_4211_im;
    _T_4213_re <= _T_4212_re;
    _T_4213_im <= _T_4212_im;
    _T_4214_re <= _T_4213_re;
    _T_4214_im <= _T_4213_im;
    _T_4215_re <= _T_4214_re;
    _T_4215_im <= _T_4214_im;
    _T_4216_re <= _T_4215_re;
    _T_4216_im <= _T_4215_im;
    _T_4217_re <= _T_4216_re;
    _T_4217_im <= _T_4216_im;
    _T_4218_re <= _T_4217_re;
    _T_4218_im <= _T_4217_im;
    _T_4219_re <= _T_4218_re;
    _T_4219_im <= _T_4218_im;
    _T_4220_re <= _T_4219_re;
    _T_4220_im <= _T_4219_im;
    _T_4221_re <= _T_4220_re;
    _T_4221_im <= _T_4220_im;
    _T_4222_re <= _T_4221_re;
    _T_4222_im <= _T_4221_im;
    _T_4223_re <= _T_4222_re;
    _T_4223_im <= _T_4222_im;
    _T_4224_re <= _T_4223_re;
    _T_4224_im <= _T_4223_im;
    _T_4225_re <= _T_4224_re;
    _T_4225_im <= _T_4224_im;
    _T_4226_re <= _T_4225_re;
    _T_4226_im <= _T_4225_im;
    _T_4227_re <= _T_4226_re;
    _T_4227_im <= _T_4226_im;
    _T_4228_re <= _T_4227_re;
    _T_4228_im <= _T_4227_im;
    _T_4229_re <= _T_4228_re;
    _T_4229_im <= _T_4228_im;
    _T_4230_re <= _T_4229_re;
    _T_4230_im <= _T_4229_im;
    _T_4231_re <= _T_4230_re;
    _T_4231_im <= _T_4230_im;
    _T_4232_re <= _T_4231_re;
    _T_4232_im <= _T_4231_im;
    _T_4233_re <= _T_4232_re;
    _T_4233_im <= _T_4232_im;
    _T_4234_re <= _T_4233_re;
    _T_4234_im <= _T_4233_im;
    _T_4235_re <= _T_4234_re;
    _T_4235_im <= _T_4234_im;
    _T_4236_re <= _T_4235_re;
    _T_4236_im <= _T_4235_im;
    _T_4237_re <= _T_4236_re;
    _T_4237_im <= _T_4236_im;
    _T_4238_re <= _T_4237_re;
    _T_4238_im <= _T_4237_im;
    _T_4239_re <= _T_4238_re;
    _T_4239_im <= _T_4238_im;
    _T_4240_re <= _T_4239_re;
    _T_4240_im <= _T_4239_im;
    _T_4241_re <= _T_4240_re;
    _T_4241_im <= _T_4240_im;
    _T_4242_re <= _T_4241_re;
    _T_4242_im <= _T_4241_im;
    _T_4243_re <= _T_4242_re;
    _T_4243_im <= _T_4242_im;
    _T_4244_re <= _T_4243_re;
    _T_4244_im <= _T_4243_im;
    _T_4245_re <= _T_4244_re;
    _T_4245_im <= _T_4244_im;
    _T_4246_re <= _T_4245_re;
    _T_4246_im <= _T_4245_im;
    _T_4247_re <= _T_4246_re;
    _T_4247_im <= _T_4246_im;
    _T_4248_re <= _T_4247_re;
    _T_4248_im <= _T_4247_im;
    _T_4249_re <= _T_4248_re;
    _T_4249_im <= _T_4248_im;
    _T_4250_re <= _T_4249_re;
    _T_4250_im <= _T_4249_im;
    _T_4251_re <= _T_4250_re;
    _T_4251_im <= _T_4250_im;
    _T_4252_re <= _T_4251_re;
    _T_4252_im <= _T_4251_im;
    _T_4253_re <= _T_4252_re;
    _T_4253_im <= _T_4252_im;
    _T_4254_re <= _T_4253_re;
    _T_4254_im <= _T_4253_im;
    _T_4255_re <= _T_4254_re;
    _T_4255_im <= _T_4254_im;
    _T_4256_re <= _T_4255_re;
    _T_4256_im <= _T_4255_im;
    _T_4257_re <= _T_4256_re;
    _T_4257_im <= _T_4256_im;
    _T_4258_re <= _T_4257_re;
    _T_4258_im <= _T_4257_im;
    _T_4259_re <= _T_4258_re;
    _T_4259_im <= _T_4258_im;
    _T_4260_re <= _T_4259_re;
    _T_4260_im <= _T_4259_im;
    _T_4261_re <= _T_4260_re;
    _T_4261_im <= _T_4260_im;
    _T_4262_re <= _T_4261_re;
    _T_4262_im <= _T_4261_im;
    _T_4263_re <= _T_4262_re;
    _T_4263_im <= _T_4262_im;
    _T_4264_re <= _T_4263_re;
    _T_4264_im <= _T_4263_im;
    _T_4265_re <= _T_4264_re;
    _T_4265_im <= _T_4264_im;
    _T_4266_re <= _T_4265_re;
    _T_4266_im <= _T_4265_im;
    _T_4267_re <= _T_4266_re;
    _T_4267_im <= _T_4266_im;
    _T_4268_re <= _T_4267_re;
    _T_4268_im <= _T_4267_im;
    _T_4269_re <= _T_4268_re;
    _T_4269_im <= _T_4268_im;
    _T_4270_re <= _T_4269_re;
    _T_4270_im <= _T_4269_im;
    _T_4271_re <= _T_4270_re;
    _T_4271_im <= _T_4270_im;
    _T_4272_re <= _T_4271_re;
    _T_4272_im <= _T_4271_im;
    _T_4273_re <= _T_4272_re;
    _T_4273_im <= _T_4272_im;
    _T_4274_re <= _T_4273_re;
    _T_4274_im <= _T_4273_im;
    _T_4275_re <= _T_4274_re;
    _T_4275_im <= _T_4274_im;
    _T_4276_re <= _T_4275_re;
    _T_4276_im <= _T_4275_im;
    _T_4277_re <= _T_4276_re;
    _T_4277_im <= _T_4276_im;
    _T_4278_re <= _T_4277_re;
    _T_4278_im <= _T_4277_im;
    _T_4279_re <= _T_4278_re;
    _T_4279_im <= _T_4278_im;
    _T_4280_re <= _T_4279_re;
    _T_4280_im <= _T_4279_im;
    _T_4281_re <= _T_4280_re;
    _T_4281_im <= _T_4280_im;
    _T_4282_re <= _T_4281_re;
    _T_4282_im <= _T_4281_im;
    _T_4283_re <= _T_4282_re;
    _T_4283_im <= _T_4282_im;
    _T_4284_re <= _T_4283_re;
    _T_4284_im <= _T_4283_im;
    _T_4285_re <= _T_4284_re;
    _T_4285_im <= _T_4284_im;
    _T_4286_re <= _T_4285_re;
    _T_4286_im <= _T_4285_im;
    _T_4287_re <= _T_4286_re;
    _T_4287_im <= _T_4286_im;
    _T_4288_re <= _T_4287_re;
    _T_4288_im <= _T_4287_im;
    _T_4289_re <= _T_4288_re;
    _T_4289_im <= _T_4288_im;
    _T_4290_re <= _T_4289_re;
    _T_4290_im <= _T_4289_im;
    _T_4291_re <= _T_4290_re;
    _T_4291_im <= _T_4290_im;
    _T_4294_re <= Butterfly_1_io_out2_re;
    _T_4294_im <= Butterfly_1_io_out2_im;
    _T_4295_re <= _T_4294_re;
    _T_4295_im <= _T_4294_im;
    _T_4296_re <= _T_4295_re;
    _T_4296_im <= _T_4295_im;
    _T_4297_re <= _T_4296_re;
    _T_4297_im <= _T_4296_im;
    _T_4298_re <= _T_4297_re;
    _T_4298_im <= _T_4297_im;
    _T_4299_re <= _T_4298_re;
    _T_4299_im <= _T_4298_im;
    _T_4300_re <= _T_4299_re;
    _T_4300_im <= _T_4299_im;
    _T_4301_re <= _T_4300_re;
    _T_4301_im <= _T_4300_im;
    _T_4302_re <= _T_4301_re;
    _T_4302_im <= _T_4301_im;
    _T_4303_re <= _T_4302_re;
    _T_4303_im <= _T_4302_im;
    _T_4304_re <= _T_4303_re;
    _T_4304_im <= _T_4303_im;
    _T_4305_re <= _T_4304_re;
    _T_4305_im <= _T_4304_im;
    _T_4306_re <= _T_4305_re;
    _T_4306_im <= _T_4305_im;
    _T_4307_re <= _T_4306_re;
    _T_4307_im <= _T_4306_im;
    _T_4308_re <= _T_4307_re;
    _T_4308_im <= _T_4307_im;
    _T_4309_re <= _T_4308_re;
    _T_4309_im <= _T_4308_im;
    _T_4310_re <= _T_4309_re;
    _T_4310_im <= _T_4309_im;
    _T_4311_re <= _T_4310_re;
    _T_4311_im <= _T_4310_im;
    _T_4312_re <= _T_4311_re;
    _T_4312_im <= _T_4311_im;
    _T_4313_re <= _T_4312_re;
    _T_4313_im <= _T_4312_im;
    _T_4314_re <= _T_4313_re;
    _T_4314_im <= _T_4313_im;
    _T_4315_re <= _T_4314_re;
    _T_4315_im <= _T_4314_im;
    _T_4316_re <= _T_4315_re;
    _T_4316_im <= _T_4315_im;
    _T_4317_re <= _T_4316_re;
    _T_4317_im <= _T_4316_im;
    _T_4318_re <= _T_4317_re;
    _T_4318_im <= _T_4317_im;
    _T_4319_re <= _T_4318_re;
    _T_4319_im <= _T_4318_im;
    _T_4320_re <= _T_4319_re;
    _T_4320_im <= _T_4319_im;
    _T_4321_re <= _T_4320_re;
    _T_4321_im <= _T_4320_im;
    _T_4322_re <= _T_4321_re;
    _T_4322_im <= _T_4321_im;
    _T_4323_re <= _T_4322_re;
    _T_4323_im <= _T_4322_im;
    _T_4324_re <= _T_4323_re;
    _T_4324_im <= _T_4323_im;
    _T_4325_re <= _T_4324_re;
    _T_4325_im <= _T_4324_im;
    _T_4326_re <= _T_4325_re;
    _T_4326_im <= _T_4325_im;
    _T_4327_re <= _T_4326_re;
    _T_4327_im <= _T_4326_im;
    _T_4328_re <= _T_4327_re;
    _T_4328_im <= _T_4327_im;
    _T_4329_re <= _T_4328_re;
    _T_4329_im <= _T_4328_im;
    _T_4330_re <= _T_4329_re;
    _T_4330_im <= _T_4329_im;
    _T_4331_re <= _T_4330_re;
    _T_4331_im <= _T_4330_im;
    _T_4332_re <= _T_4331_re;
    _T_4332_im <= _T_4331_im;
    _T_4333_re <= _T_4332_re;
    _T_4333_im <= _T_4332_im;
    _T_4334_re <= _T_4333_re;
    _T_4334_im <= _T_4333_im;
    _T_4335_re <= _T_4334_re;
    _T_4335_im <= _T_4334_im;
    _T_4336_re <= _T_4335_re;
    _T_4336_im <= _T_4335_im;
    _T_4337_re <= _T_4336_re;
    _T_4337_im <= _T_4336_im;
    _T_4338_re <= _T_4337_re;
    _T_4338_im <= _T_4337_im;
    _T_4339_re <= _T_4338_re;
    _T_4339_im <= _T_4338_im;
    _T_4340_re <= _T_4339_re;
    _T_4340_im <= _T_4339_im;
    _T_4341_re <= _T_4340_re;
    _T_4341_im <= _T_4340_im;
    _T_4342_re <= _T_4341_re;
    _T_4342_im <= _T_4341_im;
    _T_4343_re <= _T_4342_re;
    _T_4343_im <= _T_4342_im;
    _T_4344_re <= _T_4343_re;
    _T_4344_im <= _T_4343_im;
    _T_4345_re <= _T_4344_re;
    _T_4345_im <= _T_4344_im;
    _T_4346_re <= _T_4345_re;
    _T_4346_im <= _T_4345_im;
    _T_4347_re <= _T_4346_re;
    _T_4347_im <= _T_4346_im;
    _T_4348_re <= _T_4347_re;
    _T_4348_im <= _T_4347_im;
    _T_4349_re <= _T_4348_re;
    _T_4349_im <= _T_4348_im;
    _T_4350_re <= _T_4349_re;
    _T_4350_im <= _T_4349_im;
    _T_4351_re <= _T_4350_re;
    _T_4351_im <= _T_4350_im;
    _T_4352_re <= _T_4351_re;
    _T_4352_im <= _T_4351_im;
    _T_4353_re <= _T_4352_re;
    _T_4353_im <= _T_4352_im;
    _T_4354_re <= _T_4353_re;
    _T_4354_im <= _T_4353_im;
    _T_4355_re <= _T_4354_re;
    _T_4355_im <= _T_4354_im;
    _T_4356_re <= _T_4355_re;
    _T_4356_im <= _T_4355_im;
    _T_4357_re <= _T_4356_re;
    _T_4357_im <= _T_4356_im;
    _T_4358_re <= _T_4357_re;
    _T_4358_im <= _T_4357_im;
    _T_4359_re <= _T_4358_re;
    _T_4359_im <= _T_4358_im;
    _T_4360_re <= _T_4359_re;
    _T_4360_im <= _T_4359_im;
    _T_4361_re <= _T_4360_re;
    _T_4361_im <= _T_4360_im;
    _T_4362_re <= _T_4361_re;
    _T_4362_im <= _T_4361_im;
    _T_4363_re <= _T_4362_re;
    _T_4363_im <= _T_4362_im;
    _T_4364_re <= _T_4363_re;
    _T_4364_im <= _T_4363_im;
    _T_4365_re <= _T_4364_re;
    _T_4365_im <= _T_4364_im;
    _T_4366_re <= _T_4365_re;
    _T_4366_im <= _T_4365_im;
    _T_4367_re <= _T_4366_re;
    _T_4367_im <= _T_4366_im;
    _T_4368_re <= _T_4367_re;
    _T_4368_im <= _T_4367_im;
    _T_4369_re <= _T_4368_re;
    _T_4369_im <= _T_4368_im;
    _T_4370_re <= _T_4369_re;
    _T_4370_im <= _T_4369_im;
    _T_4371_re <= _T_4370_re;
    _T_4371_im <= _T_4370_im;
    _T_4372_re <= _T_4371_re;
    _T_4372_im <= _T_4371_im;
    _T_4373_re <= _T_4372_re;
    _T_4373_im <= _T_4372_im;
    _T_4374_re <= _T_4373_re;
    _T_4374_im <= _T_4373_im;
    _T_4375_re <= _T_4374_re;
    _T_4375_im <= _T_4374_im;
    _T_4376_re <= _T_4375_re;
    _T_4376_im <= _T_4375_im;
    _T_4377_re <= _T_4376_re;
    _T_4377_im <= _T_4376_im;
    _T_4378_re <= _T_4377_re;
    _T_4378_im <= _T_4377_im;
    _T_4379_re <= _T_4378_re;
    _T_4379_im <= _T_4378_im;
    _T_4380_re <= _T_4379_re;
    _T_4380_im <= _T_4379_im;
    _T_4381_re <= _T_4380_re;
    _T_4381_im <= _T_4380_im;
    _T_4382_re <= _T_4381_re;
    _T_4382_im <= _T_4381_im;
    _T_4383_re <= _T_4382_re;
    _T_4383_im <= _T_4382_im;
    _T_4384_re <= _T_4383_re;
    _T_4384_im <= _T_4383_im;
    _T_4385_re <= _T_4384_re;
    _T_4385_im <= _T_4384_im;
    _T_4386_re <= _T_4385_re;
    _T_4386_im <= _T_4385_im;
    _T_4387_re <= _T_4386_re;
    _T_4387_im <= _T_4386_im;
    _T_4388_re <= _T_4387_re;
    _T_4388_im <= _T_4387_im;
    _T_4389_re <= _T_4388_re;
    _T_4389_im <= _T_4388_im;
    _T_4390_re <= _T_4389_re;
    _T_4390_im <= _T_4389_im;
    _T_4391_re <= _T_4390_re;
    _T_4391_im <= _T_4390_im;
    _T_4392_re <= _T_4391_re;
    _T_4392_im <= _T_4391_im;
    _T_4393_re <= _T_4392_re;
    _T_4393_im <= _T_4392_im;
    _T_4394_re <= _T_4393_re;
    _T_4394_im <= _T_4393_im;
    _T_4395_re <= _T_4394_re;
    _T_4395_im <= _T_4394_im;
    _T_4396_re <= _T_4395_re;
    _T_4396_im <= _T_4395_im;
    _T_4397_re <= _T_4396_re;
    _T_4397_im <= _T_4396_im;
    _T_4398_re <= _T_4397_re;
    _T_4398_im <= _T_4397_im;
    _T_4399_re <= _T_4398_re;
    _T_4399_im <= _T_4398_im;
    _T_4400_re <= _T_4399_re;
    _T_4400_im <= _T_4399_im;
    _T_4401_re <= _T_4400_re;
    _T_4401_im <= _T_4400_im;
    _T_4402_re <= _T_4401_re;
    _T_4402_im <= _T_4401_im;
    _T_4403_re <= _T_4402_re;
    _T_4403_im <= _T_4402_im;
    _T_4404_re <= _T_4403_re;
    _T_4404_im <= _T_4403_im;
    _T_4405_re <= _T_4404_re;
    _T_4405_im <= _T_4404_im;
    _T_4406_re <= _T_4405_re;
    _T_4406_im <= _T_4405_im;
    _T_4407_re <= _T_4406_re;
    _T_4407_im <= _T_4406_im;
    _T_4408_re <= _T_4407_re;
    _T_4408_im <= _T_4407_im;
    _T_4409_re <= _T_4408_re;
    _T_4409_im <= _T_4408_im;
    _T_4410_re <= _T_4409_re;
    _T_4410_im <= _T_4409_im;
    _T_4411_re <= _T_4410_re;
    _T_4411_im <= _T_4410_im;
    _T_4412_re <= _T_4411_re;
    _T_4412_im <= _T_4411_im;
    _T_4413_re <= _T_4412_re;
    _T_4413_im <= _T_4412_im;
    _T_4414_re <= _T_4413_re;
    _T_4414_im <= _T_4413_im;
    _T_4415_re <= _T_4414_re;
    _T_4415_im <= _T_4414_im;
    _T_4416_re <= _T_4415_re;
    _T_4416_im <= _T_4415_im;
    _T_4417_re <= _T_4416_re;
    _T_4417_im <= _T_4416_im;
    _T_4418_re <= _T_4417_re;
    _T_4418_im <= _T_4417_im;
    _T_4419_re <= _T_4418_re;
    _T_4419_im <= _T_4418_im;
    _T_4420_re <= _T_4419_re;
    _T_4420_im <= _T_4419_im;
    _T_4421_re <= _T_4420_re;
    _T_4421_im <= _T_4420_im;
    _T_4422_re <= _T_4421_re;
    _T_4422_im <= _T_4421_im;
    _T_4423_re <= _T_4422_re;
    _T_4423_im <= _T_4422_im;
    _T_4424_re <= _T_4423_re;
    _T_4424_im <= _T_4423_im;
    _T_4425_re <= _T_4424_re;
    _T_4425_im <= _T_4424_im;
    _T_4426_re <= _T_4425_re;
    _T_4426_im <= _T_4425_im;
    _T_4427_re <= _T_4426_re;
    _T_4427_im <= _T_4426_im;
    _T_4428_re <= _T_4427_re;
    _T_4428_im <= _T_4427_im;
    _T_4429_re <= _T_4428_re;
    _T_4429_im <= _T_4428_im;
    _T_4430_re <= _T_4429_re;
    _T_4430_im <= _T_4429_im;
    _T_4431_re <= _T_4430_re;
    _T_4431_im <= _T_4430_im;
    _T_4432_re <= _T_4431_re;
    _T_4432_im <= _T_4431_im;
    _T_4433_re <= _T_4432_re;
    _T_4433_im <= _T_4432_im;
    _T_4434_re <= _T_4433_re;
    _T_4434_im <= _T_4433_im;
    _T_4435_re <= _T_4434_re;
    _T_4435_im <= _T_4434_im;
    _T_4436_re <= _T_4435_re;
    _T_4436_im <= _T_4435_im;
    _T_4437_re <= _T_4436_re;
    _T_4437_im <= _T_4436_im;
    _T_4438_re <= _T_4437_re;
    _T_4438_im <= _T_4437_im;
    _T_4439_re <= _T_4438_re;
    _T_4439_im <= _T_4438_im;
    _T_4440_re <= _T_4439_re;
    _T_4440_im <= _T_4439_im;
    _T_4441_re <= _T_4440_re;
    _T_4441_im <= _T_4440_im;
    _T_4442_re <= _T_4441_re;
    _T_4442_im <= _T_4441_im;
    _T_4443_re <= _T_4442_re;
    _T_4443_im <= _T_4442_im;
    _T_4444_re <= _T_4443_re;
    _T_4444_im <= _T_4443_im;
    _T_4445_re <= _T_4444_re;
    _T_4445_im <= _T_4444_im;
    _T_4446_re <= _T_4445_re;
    _T_4446_im <= _T_4445_im;
    _T_4447_re <= _T_4446_re;
    _T_4447_im <= _T_4446_im;
    _T_4448_re <= _T_4447_re;
    _T_4448_im <= _T_4447_im;
    _T_4449_re <= _T_4448_re;
    _T_4449_im <= _T_4448_im;
    _T_4450_re <= _T_4449_re;
    _T_4450_im <= _T_4449_im;
    _T_4451_re <= _T_4450_re;
    _T_4451_im <= _T_4450_im;
    _T_4452_re <= _T_4451_re;
    _T_4452_im <= _T_4451_im;
    _T_4453_re <= _T_4452_re;
    _T_4453_im <= _T_4452_im;
    _T_4454_re <= _T_4453_re;
    _T_4454_im <= _T_4453_im;
    _T_4455_re <= _T_4454_re;
    _T_4455_im <= _T_4454_im;
    _T_4456_re <= _T_4455_re;
    _T_4456_im <= _T_4455_im;
    _T_4457_re <= _T_4456_re;
    _T_4457_im <= _T_4456_im;
    _T_4458_re <= _T_4457_re;
    _T_4458_im <= _T_4457_im;
    _T_4459_re <= _T_4458_re;
    _T_4459_im <= _T_4458_im;
    _T_4460_re <= _T_4459_re;
    _T_4460_im <= _T_4459_im;
    _T_4461_re <= _T_4460_re;
    _T_4461_im <= _T_4460_im;
    _T_4462_re <= _T_4461_re;
    _T_4462_im <= _T_4461_im;
    _T_4463_re <= _T_4462_re;
    _T_4463_im <= _T_4462_im;
    _T_4464_re <= _T_4463_re;
    _T_4464_im <= _T_4463_im;
    _T_4465_re <= _T_4464_re;
    _T_4465_im <= _T_4464_im;
    _T_4466_re <= _T_4465_re;
    _T_4466_im <= _T_4465_im;
    _T_4467_re <= _T_4466_re;
    _T_4467_im <= _T_4466_im;
    _T_4468_re <= _T_4467_re;
    _T_4468_im <= _T_4467_im;
    _T_4469_re <= _T_4468_re;
    _T_4469_im <= _T_4468_im;
    _T_4470_re <= _T_4469_re;
    _T_4470_im <= _T_4469_im;
    _T_4471_re <= _T_4470_re;
    _T_4471_im <= _T_4470_im;
    _T_4472_re <= _T_4471_re;
    _T_4472_im <= _T_4471_im;
    _T_4473_re <= _T_4472_re;
    _T_4473_im <= _T_4472_im;
    _T_4474_re <= _T_4473_re;
    _T_4474_im <= _T_4473_im;
    _T_4475_re <= _T_4474_re;
    _T_4475_im <= _T_4474_im;
    _T_4476_re <= _T_4475_re;
    _T_4476_im <= _T_4475_im;
    _T_4477_re <= _T_4476_re;
    _T_4477_im <= _T_4476_im;
    _T_4478_re <= _T_4477_re;
    _T_4478_im <= _T_4477_im;
    _T_4479_re <= _T_4478_re;
    _T_4479_im <= _T_4478_im;
    _T_4480_re <= _T_4479_re;
    _T_4480_im <= _T_4479_im;
    _T_4481_re <= _T_4480_re;
    _T_4481_im <= _T_4480_im;
    _T_4482_re <= _T_4481_re;
    _T_4482_im <= _T_4481_im;
    _T_4483_re <= _T_4482_re;
    _T_4483_im <= _T_4482_im;
    _T_4484_re <= _T_4483_re;
    _T_4484_im <= _T_4483_im;
    _T_4485_re <= _T_4484_re;
    _T_4485_im <= _T_4484_im;
    _T_4486_re <= _T_4485_re;
    _T_4486_im <= _T_4485_im;
    _T_4487_re <= _T_4486_re;
    _T_4487_im <= _T_4486_im;
    _T_4488_re <= _T_4487_re;
    _T_4488_im <= _T_4487_im;
    _T_4489_re <= _T_4488_re;
    _T_4489_im <= _T_4488_im;
    _T_4490_re <= _T_4489_re;
    _T_4490_im <= _T_4489_im;
    _T_4491_re <= _T_4490_re;
    _T_4491_im <= _T_4490_im;
    _T_4492_re <= _T_4491_re;
    _T_4492_im <= _T_4491_im;
    _T_4493_re <= _T_4492_re;
    _T_4493_im <= _T_4492_im;
    _T_4494_re <= _T_4493_re;
    _T_4494_im <= _T_4493_im;
    _T_4495_re <= _T_4494_re;
    _T_4495_im <= _T_4494_im;
    _T_4496_re <= _T_4495_re;
    _T_4496_im <= _T_4495_im;
    _T_4497_re <= _T_4496_re;
    _T_4497_im <= _T_4496_im;
    _T_4498_re <= _T_4497_re;
    _T_4498_im <= _T_4497_im;
    _T_4499_re <= _T_4498_re;
    _T_4499_im <= _T_4498_im;
    _T_4500_re <= _T_4499_re;
    _T_4500_im <= _T_4499_im;
    _T_4501_re <= _T_4500_re;
    _T_4501_im <= _T_4500_im;
    _T_4502_re <= _T_4501_re;
    _T_4502_im <= _T_4501_im;
    _T_4503_re <= _T_4502_re;
    _T_4503_im <= _T_4502_im;
    _T_4504_re <= _T_4503_re;
    _T_4504_im <= _T_4503_im;
    _T_4505_re <= _T_4504_re;
    _T_4505_im <= _T_4504_im;
    _T_4506_re <= _T_4505_re;
    _T_4506_im <= _T_4505_im;
    _T_4507_re <= _T_4506_re;
    _T_4507_im <= _T_4506_im;
    _T_4508_re <= _T_4507_re;
    _T_4508_im <= _T_4507_im;
    _T_4509_re <= _T_4508_re;
    _T_4509_im <= _T_4508_im;
    _T_4510_re <= _T_4509_re;
    _T_4510_im <= _T_4509_im;
    _T_4511_re <= _T_4510_re;
    _T_4511_im <= _T_4510_im;
    _T_4512_re <= _T_4511_re;
    _T_4512_im <= _T_4511_im;
    _T_4513_re <= _T_4512_re;
    _T_4513_im <= _T_4512_im;
    _T_4514_re <= _T_4513_re;
    _T_4514_im <= _T_4513_im;
    _T_4515_re <= _T_4514_re;
    _T_4515_im <= _T_4514_im;
    _T_4516_re <= _T_4515_re;
    _T_4516_im <= _T_4515_im;
    _T_4517_re <= _T_4516_re;
    _T_4517_im <= _T_4516_im;
    _T_4518_re <= _T_4517_re;
    _T_4518_im <= _T_4517_im;
    _T_4519_re <= _T_4518_re;
    _T_4519_im <= _T_4518_im;
    _T_4520_re <= _T_4519_re;
    _T_4520_im <= _T_4519_im;
    _T_4521_re <= _T_4520_re;
    _T_4521_im <= _T_4520_im;
    _T_4522_re <= _T_4521_re;
    _T_4522_im <= _T_4521_im;
    _T_4523_re <= _T_4522_re;
    _T_4523_im <= _T_4522_im;
    _T_4524_re <= _T_4523_re;
    _T_4524_im <= _T_4523_im;
    _T_4525_re <= _T_4524_re;
    _T_4525_im <= _T_4524_im;
    _T_4526_re <= _T_4525_re;
    _T_4526_im <= _T_4525_im;
    _T_4527_re <= _T_4526_re;
    _T_4527_im <= _T_4526_im;
    _T_4528_re <= _T_4527_re;
    _T_4528_im <= _T_4527_im;
    _T_4529_re <= _T_4528_re;
    _T_4529_im <= _T_4528_im;
    _T_4530_re <= _T_4529_re;
    _T_4530_im <= _T_4529_im;
    _T_4531_re <= _T_4530_re;
    _T_4531_im <= _T_4530_im;
    _T_4532_re <= _T_4531_re;
    _T_4532_im <= _T_4531_im;
    _T_4533_re <= _T_4532_re;
    _T_4533_im <= _T_4532_im;
    _T_4534_re <= _T_4533_re;
    _T_4534_im <= _T_4533_im;
    _T_4535_re <= _T_4534_re;
    _T_4535_im <= _T_4534_im;
    _T_4536_re <= _T_4535_re;
    _T_4536_im <= _T_4535_im;
    _T_4537_re <= _T_4536_re;
    _T_4537_im <= _T_4536_im;
    _T_4538_re <= _T_4537_re;
    _T_4538_im <= _T_4537_im;
    _T_4539_re <= _T_4538_re;
    _T_4539_im <= _T_4538_im;
    _T_4540_re <= _T_4539_re;
    _T_4540_im <= _T_4539_im;
    _T_4541_re <= _T_4540_re;
    _T_4541_im <= _T_4540_im;
    _T_4542_re <= _T_4541_re;
    _T_4542_im <= _T_4541_im;
    _T_4543_re <= _T_4542_re;
    _T_4543_im <= _T_4542_im;
    _T_4544_re <= _T_4543_re;
    _T_4544_im <= _T_4543_im;
    _T_4545_re <= _T_4544_re;
    _T_4545_im <= _T_4544_im;
    _T_4546_re <= _T_4545_re;
    _T_4546_im <= _T_4545_im;
    _T_4547_re <= _T_4546_re;
    _T_4547_im <= _T_4546_im;
    _T_4548_re <= _T_4547_re;
    _T_4548_im <= _T_4547_im;
    _T_4549_re <= _T_4548_re;
    _T_4549_im <= _T_4548_im;
    _T_4550_re <= _T_4549_re;
    _T_4550_im <= _T_4549_im;
    _T_4551_re <= _T_4550_re;
    _T_4551_im <= _T_4550_im;
    _T_4552_re <= _T_4551_re;
    _T_4552_im <= _T_4551_im;
    _T_4553_re <= _T_4552_re;
    _T_4553_im <= _T_4552_im;
    _T_4554_re <= _T_4553_re;
    _T_4554_im <= _T_4553_im;
    _T_4555_re <= _T_4554_re;
    _T_4555_im <= _T_4554_im;
    _T_4556_re <= _T_4555_re;
    _T_4556_im <= _T_4555_im;
    _T_4557_re <= _T_4556_re;
    _T_4557_im <= _T_4556_im;
    _T_4558_re <= _T_4557_re;
    _T_4558_im <= _T_4557_im;
    _T_4559_re <= _T_4558_re;
    _T_4559_im <= _T_4558_im;
    _T_4560_re <= _T_4559_re;
    _T_4560_im <= _T_4559_im;
    _T_4561_re <= _T_4560_re;
    _T_4561_im <= _T_4560_im;
    _T_4562_re <= _T_4561_re;
    _T_4562_im <= _T_4561_im;
    _T_4563_re <= _T_4562_re;
    _T_4563_im <= _T_4562_im;
    _T_4564_re <= _T_4563_re;
    _T_4564_im <= _T_4563_im;
    _T_4565_re <= _T_4564_re;
    _T_4565_im <= _T_4564_im;
    _T_4566_re <= _T_4565_re;
    _T_4566_im <= _T_4565_im;
    _T_4567_re <= _T_4566_re;
    _T_4567_im <= _T_4566_im;
    _T_4568_re <= _T_4567_re;
    _T_4568_im <= _T_4567_im;
    _T_4569_re <= _T_4568_re;
    _T_4569_im <= _T_4568_im;
    _T_4570_re <= _T_4569_re;
    _T_4570_im <= _T_4569_im;
    _T_4571_re <= _T_4570_re;
    _T_4571_im <= _T_4570_im;
    _T_4572_re <= _T_4571_re;
    _T_4572_im <= _T_4571_im;
    _T_4573_re <= _T_4572_re;
    _T_4573_im <= _T_4572_im;
    _T_4574_re <= _T_4573_re;
    _T_4574_im <= _T_4573_im;
    _T_4575_re <= _T_4574_re;
    _T_4575_im <= _T_4574_im;
    _T_4576_re <= _T_4575_re;
    _T_4576_im <= _T_4575_im;
    _T_4577_re <= _T_4576_re;
    _T_4577_im <= _T_4576_im;
    _T_4578_re <= _T_4577_re;
    _T_4578_im <= _T_4577_im;
    _T_4579_re <= _T_4578_re;
    _T_4579_im <= _T_4578_im;
    _T_4580_re <= _T_4579_re;
    _T_4580_im <= _T_4579_im;
    _T_4581_re <= _T_4580_re;
    _T_4581_im <= _T_4580_im;
    _T_4582_re <= _T_4581_re;
    _T_4582_im <= _T_4581_im;
    _T_4583_re <= _T_4582_re;
    _T_4583_im <= _T_4582_im;
    _T_4584_re <= _T_4583_re;
    _T_4584_im <= _T_4583_im;
    _T_4585_re <= _T_4584_re;
    _T_4585_im <= _T_4584_im;
    _T_4586_re <= _T_4585_re;
    _T_4586_im <= _T_4585_im;
    _T_4587_re <= _T_4586_re;
    _T_4587_im <= _T_4586_im;
    _T_4588_re <= _T_4587_re;
    _T_4588_im <= _T_4587_im;
    _T_4589_re <= _T_4588_re;
    _T_4589_im <= _T_4588_im;
    _T_4590_re <= _T_4589_re;
    _T_4590_im <= _T_4589_im;
    _T_4591_re <= _T_4590_re;
    _T_4591_im <= _T_4590_im;
    _T_4592_re <= _T_4591_re;
    _T_4592_im <= _T_4591_im;
    _T_4593_re <= _T_4592_re;
    _T_4593_im <= _T_4592_im;
    _T_4594_re <= _T_4593_re;
    _T_4594_im <= _T_4593_im;
    _T_4595_re <= _T_4594_re;
    _T_4595_im <= _T_4594_im;
    _T_4596_re <= _T_4595_re;
    _T_4596_im <= _T_4595_im;
    _T_4597_re <= _T_4596_re;
    _T_4597_im <= _T_4596_im;
    _T_4598_re <= _T_4597_re;
    _T_4598_im <= _T_4597_im;
    _T_4599_re <= _T_4598_re;
    _T_4599_im <= _T_4598_im;
    _T_4600_re <= _T_4599_re;
    _T_4600_im <= _T_4599_im;
    _T_4601_re <= _T_4600_re;
    _T_4601_im <= _T_4600_im;
    _T_4602_re <= _T_4601_re;
    _T_4602_im <= _T_4601_im;
    _T_4603_re <= _T_4602_re;
    _T_4603_im <= _T_4602_im;
    _T_4604_re <= _T_4603_re;
    _T_4604_im <= _T_4603_im;
    _T_4605_re <= _T_4604_re;
    _T_4605_im <= _T_4604_im;
    _T_4606_re <= _T_4605_re;
    _T_4606_im <= _T_4605_im;
    _T_4607_re <= _T_4606_re;
    _T_4607_im <= _T_4606_im;
    _T_4608_re <= _T_4607_re;
    _T_4608_im <= _T_4607_im;
    _T_4609_re <= _T_4608_re;
    _T_4609_im <= _T_4608_im;
    _T_4610_re <= _T_4609_re;
    _T_4610_im <= _T_4609_im;
    _T_4611_re <= _T_4610_re;
    _T_4611_im <= _T_4610_im;
    _T_4612_re <= _T_4611_re;
    _T_4612_im <= _T_4611_im;
    _T_4613_re <= _T_4612_re;
    _T_4613_im <= _T_4612_im;
    _T_4614_re <= _T_4613_re;
    _T_4614_im <= _T_4613_im;
    _T_4615_re <= _T_4614_re;
    _T_4615_im <= _T_4614_im;
    _T_4616_re <= _T_4615_re;
    _T_4616_im <= _T_4615_im;
    _T_4617_re <= _T_4616_re;
    _T_4617_im <= _T_4616_im;
    _T_4618_re <= _T_4617_re;
    _T_4618_im <= _T_4617_im;
    _T_4619_re <= _T_4618_re;
    _T_4619_im <= _T_4618_im;
    _T_4620_re <= _T_4619_re;
    _T_4620_im <= _T_4619_im;
    _T_4621_re <= _T_4620_re;
    _T_4621_im <= _T_4620_im;
    _T_4622_re <= _T_4621_re;
    _T_4622_im <= _T_4621_im;
    _T_4623_re <= _T_4622_re;
    _T_4623_im <= _T_4622_im;
    _T_4624_re <= _T_4623_re;
    _T_4624_im <= _T_4623_im;
    _T_4625_re <= _T_4624_re;
    _T_4625_im <= _T_4624_im;
    _T_4626_re <= _T_4625_re;
    _T_4626_im <= _T_4625_im;
    _T_4627_re <= _T_4626_re;
    _T_4627_im <= _T_4626_im;
    _T_4628_re <= _T_4627_re;
    _T_4628_im <= _T_4627_im;
    _T_4629_re <= _T_4628_re;
    _T_4629_im <= _T_4628_im;
    _T_4630_re <= _T_4629_re;
    _T_4630_im <= _T_4629_im;
    _T_4631_re <= _T_4630_re;
    _T_4631_im <= _T_4630_im;
    _T_4632_re <= _T_4631_re;
    _T_4632_im <= _T_4631_im;
    _T_4633_re <= _T_4632_re;
    _T_4633_im <= _T_4632_im;
    _T_4634_re <= _T_4633_re;
    _T_4634_im <= _T_4633_im;
    _T_4635_re <= _T_4634_re;
    _T_4635_im <= _T_4634_im;
    _T_4636_re <= _T_4635_re;
    _T_4636_im <= _T_4635_im;
    _T_4637_re <= _T_4636_re;
    _T_4637_im <= _T_4636_im;
    _T_4638_re <= _T_4637_re;
    _T_4638_im <= _T_4637_im;
    _T_4639_re <= _T_4638_re;
    _T_4639_im <= _T_4638_im;
    _T_4640_re <= _T_4639_re;
    _T_4640_im <= _T_4639_im;
    _T_4641_re <= _T_4640_re;
    _T_4641_im <= _T_4640_im;
    _T_4642_re <= _T_4641_re;
    _T_4642_im <= _T_4641_im;
    _T_4643_re <= _T_4642_re;
    _T_4643_im <= _T_4642_im;
    _T_4644_re <= _T_4643_re;
    _T_4644_im <= _T_4643_im;
    _T_4645_re <= _T_4644_re;
    _T_4645_im <= _T_4644_im;
    _T_4646_re <= _T_4645_re;
    _T_4646_im <= _T_4645_im;
    _T_4647_re <= _T_4646_re;
    _T_4647_im <= _T_4646_im;
    _T_4648_re <= _T_4647_re;
    _T_4648_im <= _T_4647_im;
    _T_4649_re <= _T_4648_re;
    _T_4649_im <= _T_4648_im;
    _T_4650_re <= _T_4649_re;
    _T_4650_im <= _T_4649_im;
    _T_4651_re <= _T_4650_re;
    _T_4651_im <= _T_4650_im;
    _T_4652_re <= _T_4651_re;
    _T_4652_im <= _T_4651_im;
    _T_4653_re <= _T_4652_re;
    _T_4653_im <= _T_4652_im;
    _T_4654_re <= _T_4653_re;
    _T_4654_im <= _T_4653_im;
    _T_4655_re <= _T_4654_re;
    _T_4655_im <= _T_4654_im;
    _T_4656_re <= _T_4655_re;
    _T_4656_im <= _T_4655_im;
    _T_4657_re <= _T_4656_re;
    _T_4657_im <= _T_4656_im;
    _T_4658_re <= _T_4657_re;
    _T_4658_im <= _T_4657_im;
    _T_4659_re <= _T_4658_re;
    _T_4659_im <= _T_4658_im;
    _T_4660_re <= _T_4659_re;
    _T_4660_im <= _T_4659_im;
    _T_4661_re <= _T_4660_re;
    _T_4661_im <= _T_4660_im;
    _T_4662_re <= _T_4661_re;
    _T_4662_im <= _T_4661_im;
    _T_4663_re <= _T_4662_re;
    _T_4663_im <= _T_4662_im;
    _T_4664_re <= _T_4663_re;
    _T_4664_im <= _T_4663_im;
    _T_4665_re <= _T_4664_re;
    _T_4665_im <= _T_4664_im;
    _T_4666_re <= _T_4665_re;
    _T_4666_im <= _T_4665_im;
    _T_4667_re <= _T_4666_re;
    _T_4667_im <= _T_4666_im;
    _T_4668_re <= _T_4667_re;
    _T_4668_im <= _T_4667_im;
    _T_4669_re <= _T_4668_re;
    _T_4669_im <= _T_4668_im;
    _T_4670_re <= _T_4669_re;
    _T_4670_im <= _T_4669_im;
    _T_4671_re <= _T_4670_re;
    _T_4671_im <= _T_4670_im;
    _T_4672_re <= _T_4671_re;
    _T_4672_im <= _T_4671_im;
    _T_4673_re <= _T_4672_re;
    _T_4673_im <= _T_4672_im;
    _T_4674_re <= _T_4673_re;
    _T_4674_im <= _T_4673_im;
    _T_4675_re <= _T_4674_re;
    _T_4675_im <= _T_4674_im;
    _T_4676_re <= _T_4675_re;
    _T_4676_im <= _T_4675_im;
    _T_4677_re <= _T_4676_re;
    _T_4677_im <= _T_4676_im;
    _T_4678_re <= _T_4677_re;
    _T_4678_im <= _T_4677_im;
    _T_4679_re <= _T_4678_re;
    _T_4679_im <= _T_4678_im;
    _T_4680_re <= _T_4679_re;
    _T_4680_im <= _T_4679_im;
    _T_4681_re <= _T_4680_re;
    _T_4681_im <= _T_4680_im;
    _T_4682_re <= _T_4681_re;
    _T_4682_im <= _T_4681_im;
    _T_4683_re <= _T_4682_re;
    _T_4683_im <= _T_4682_im;
    _T_4684_re <= _T_4683_re;
    _T_4684_im <= _T_4683_im;
    _T_4685_re <= _T_4684_re;
    _T_4685_im <= _T_4684_im;
    _T_4686_re <= _T_4685_re;
    _T_4686_im <= _T_4685_im;
    _T_4687_re <= _T_4686_re;
    _T_4687_im <= _T_4686_im;
    _T_4688_re <= _T_4687_re;
    _T_4688_im <= _T_4687_im;
    _T_4689_re <= _T_4688_re;
    _T_4689_im <= _T_4688_im;
    _T_4690_re <= _T_4689_re;
    _T_4690_im <= _T_4689_im;
    _T_4691_re <= _T_4690_re;
    _T_4691_im <= _T_4690_im;
    _T_4692_re <= _T_4691_re;
    _T_4692_im <= _T_4691_im;
    _T_4693_re <= _T_4692_re;
    _T_4693_im <= _T_4692_im;
    _T_4694_re <= _T_4693_re;
    _T_4694_im <= _T_4693_im;
    _T_4695_re <= _T_4694_re;
    _T_4695_im <= _T_4694_im;
    _T_4696_re <= _T_4695_re;
    _T_4696_im <= _T_4695_im;
    _T_4697_re <= _T_4696_re;
    _T_4697_im <= _T_4696_im;
    _T_4698_re <= _T_4697_re;
    _T_4698_im <= _T_4697_im;
    _T_4699_re <= _T_4698_re;
    _T_4699_im <= _T_4698_im;
    _T_4700_re <= _T_4699_re;
    _T_4700_im <= _T_4699_im;
    _T_4701_re <= _T_4700_re;
    _T_4701_im <= _T_4700_im;
    _T_4702_re <= _T_4701_re;
    _T_4702_im <= _T_4701_im;
    _T_4703_re <= _T_4702_re;
    _T_4703_im <= _T_4702_im;
    _T_4704_re <= _T_4703_re;
    _T_4704_im <= _T_4703_im;
    _T_4705_re <= _T_4704_re;
    _T_4705_im <= _T_4704_im;
    _T_4706_re <= _T_4705_re;
    _T_4706_im <= _T_4705_im;
    _T_4707_re <= _T_4706_re;
    _T_4707_im <= _T_4706_im;
    _T_4708_re <= _T_4707_re;
    _T_4708_im <= _T_4707_im;
    _T_4709_re <= _T_4708_re;
    _T_4709_im <= _T_4708_im;
    _T_4710_re <= _T_4709_re;
    _T_4710_im <= _T_4709_im;
    _T_4711_re <= _T_4710_re;
    _T_4711_im <= _T_4710_im;
    _T_4712_re <= _T_4711_re;
    _T_4712_im <= _T_4711_im;
    _T_4713_re <= _T_4712_re;
    _T_4713_im <= _T_4712_im;
    _T_4714_re <= _T_4713_re;
    _T_4714_im <= _T_4713_im;
    _T_4715_re <= _T_4714_re;
    _T_4715_im <= _T_4714_im;
    _T_4716_re <= _T_4715_re;
    _T_4716_im <= _T_4715_im;
    _T_4717_re <= _T_4716_re;
    _T_4717_im <= _T_4716_im;
    _T_4718_re <= _T_4717_re;
    _T_4718_im <= _T_4717_im;
    _T_4719_re <= _T_4718_re;
    _T_4719_im <= _T_4718_im;
    _T_4720_re <= _T_4719_re;
    _T_4720_im <= _T_4719_im;
    _T_4721_re <= _T_4720_re;
    _T_4721_im <= _T_4720_im;
    _T_4722_re <= _T_4721_re;
    _T_4722_im <= _T_4721_im;
    _T_4723_re <= _T_4722_re;
    _T_4723_im <= _T_4722_im;
    _T_4724_re <= _T_4723_re;
    _T_4724_im <= _T_4723_im;
    _T_4725_re <= _T_4724_re;
    _T_4725_im <= _T_4724_im;
    _T_4726_re <= _T_4725_re;
    _T_4726_im <= _T_4725_im;
    _T_4727_re <= _T_4726_re;
    _T_4727_im <= _T_4726_im;
    _T_4728_re <= _T_4727_re;
    _T_4728_im <= _T_4727_im;
    _T_4729_re <= _T_4728_re;
    _T_4729_im <= _T_4728_im;
    _T_4730_re <= _T_4729_re;
    _T_4730_im <= _T_4729_im;
    _T_4731_re <= _T_4730_re;
    _T_4731_im <= _T_4730_im;
    _T_4732_re <= _T_4731_re;
    _T_4732_im <= _T_4731_im;
    _T_4733_re <= _T_4732_re;
    _T_4733_im <= _T_4732_im;
    _T_4734_re <= _T_4733_re;
    _T_4734_im <= _T_4733_im;
    _T_4735_re <= _T_4734_re;
    _T_4735_im <= _T_4734_im;
    _T_4736_re <= _T_4735_re;
    _T_4736_im <= _T_4735_im;
    _T_4737_re <= _T_4736_re;
    _T_4737_im <= _T_4736_im;
    _T_4738_re <= _T_4737_re;
    _T_4738_im <= _T_4737_im;
    _T_4739_re <= _T_4738_re;
    _T_4739_im <= _T_4738_im;
    _T_4740_re <= _T_4739_re;
    _T_4740_im <= _T_4739_im;
    _T_4741_re <= _T_4740_re;
    _T_4741_im <= _T_4740_im;
    _T_4742_re <= _T_4741_re;
    _T_4742_im <= _T_4741_im;
    _T_4743_re <= _T_4742_re;
    _T_4743_im <= _T_4742_im;
    _T_4744_re <= _T_4743_re;
    _T_4744_im <= _T_4743_im;
    _T_4745_re <= _T_4744_re;
    _T_4745_im <= _T_4744_im;
    _T_4746_re <= _T_4745_re;
    _T_4746_im <= _T_4745_im;
    _T_4747_re <= _T_4746_re;
    _T_4747_im <= _T_4746_im;
    _T_4748_re <= _T_4747_re;
    _T_4748_im <= _T_4747_im;
    _T_4749_re <= _T_4748_re;
    _T_4749_im <= _T_4748_im;
    _T_4750_re <= _T_4749_re;
    _T_4750_im <= _T_4749_im;
    _T_4751_re <= _T_4750_re;
    _T_4751_im <= _T_4750_im;
    _T_4752_re <= _T_4751_re;
    _T_4752_im <= _T_4751_im;
    _T_4753_re <= _T_4752_re;
    _T_4753_im <= _T_4752_im;
    _T_4754_re <= _T_4753_re;
    _T_4754_im <= _T_4753_im;
    _T_4755_re <= _T_4754_re;
    _T_4755_im <= _T_4754_im;
    _T_4756_re <= _T_4755_re;
    _T_4756_im <= _T_4755_im;
    _T_4757_re <= _T_4756_re;
    _T_4757_im <= _T_4756_im;
    _T_4758_re <= _T_4757_re;
    _T_4758_im <= _T_4757_im;
    _T_4759_re <= _T_4758_re;
    _T_4759_im <= _T_4758_im;
    _T_4760_re <= _T_4759_re;
    _T_4760_im <= _T_4759_im;
    _T_4761_re <= _T_4760_re;
    _T_4761_im <= _T_4760_im;
    _T_4762_re <= _T_4761_re;
    _T_4762_im <= _T_4761_im;
    _T_4763_re <= _T_4762_re;
    _T_4763_im <= _T_4762_im;
    _T_4764_re <= _T_4763_re;
    _T_4764_im <= _T_4763_im;
    _T_4765_re <= _T_4764_re;
    _T_4765_im <= _T_4764_im;
    _T_4766_re <= _T_4765_re;
    _T_4766_im <= _T_4765_im;
    _T_4767_re <= _T_4766_re;
    _T_4767_im <= _T_4766_im;
    _T_4768_re <= _T_4767_re;
    _T_4768_im <= _T_4767_im;
    _T_4769_re <= _T_4768_re;
    _T_4769_im <= _T_4768_im;
    _T_4770_re <= _T_4769_re;
    _T_4770_im <= _T_4769_im;
    _T_4771_re <= _T_4770_re;
    _T_4771_im <= _T_4770_im;
    _T_4772_re <= _T_4771_re;
    _T_4772_im <= _T_4771_im;
    _T_4773_re <= _T_4772_re;
    _T_4773_im <= _T_4772_im;
    _T_4774_re <= _T_4773_re;
    _T_4774_im <= _T_4773_im;
    _T_4775_re <= _T_4774_re;
    _T_4775_im <= _T_4774_im;
    _T_4776_re <= _T_4775_re;
    _T_4776_im <= _T_4775_im;
    _T_4777_re <= _T_4776_re;
    _T_4777_im <= _T_4776_im;
    _T_4778_re <= _T_4777_re;
    _T_4778_im <= _T_4777_im;
    _T_4779_re <= _T_4778_re;
    _T_4779_im <= _T_4778_im;
    _T_4780_re <= _T_4779_re;
    _T_4780_im <= _T_4779_im;
    _T_4781_re <= _T_4780_re;
    _T_4781_im <= _T_4780_im;
    _T_4782_re <= _T_4781_re;
    _T_4782_im <= _T_4781_im;
    _T_4783_re <= _T_4782_re;
    _T_4783_im <= _T_4782_im;
    _T_4784_re <= _T_4783_re;
    _T_4784_im <= _T_4783_im;
    _T_4785_re <= _T_4784_re;
    _T_4785_im <= _T_4784_im;
    _T_4786_re <= _T_4785_re;
    _T_4786_im <= _T_4785_im;
    _T_4787_re <= _T_4786_re;
    _T_4787_im <= _T_4786_im;
    _T_4788_re <= _T_4787_re;
    _T_4788_im <= _T_4787_im;
    _T_4789_re <= _T_4788_re;
    _T_4789_im <= _T_4788_im;
    _T_4790_re <= _T_4789_re;
    _T_4790_im <= _T_4789_im;
    _T_4791_re <= _T_4790_re;
    _T_4791_im <= _T_4790_im;
    _T_4792_re <= _T_4791_re;
    _T_4792_im <= _T_4791_im;
    _T_4793_re <= _T_4792_re;
    _T_4793_im <= _T_4792_im;
    _T_4794_re <= _T_4793_re;
    _T_4794_im <= _T_4793_im;
    _T_4795_re <= _T_4794_re;
    _T_4795_im <= _T_4794_im;
    _T_4796_re <= _T_4795_re;
    _T_4796_im <= _T_4795_im;
    _T_4797_re <= _T_4796_re;
    _T_4797_im <= _T_4796_im;
    _T_4798_re <= _T_4797_re;
    _T_4798_im <= _T_4797_im;
    _T_4799_re <= _T_4798_re;
    _T_4799_im <= _T_4798_im;
    _T_4800_re <= _T_4799_re;
    _T_4800_im <= _T_4799_im;
    _T_4801_re <= _T_4800_re;
    _T_4801_im <= _T_4800_im;
    _T_4802_re <= _T_4801_re;
    _T_4802_im <= _T_4801_im;
    _T_4803_re <= _T_4802_re;
    _T_4803_im <= _T_4802_im;
    _T_4804_re <= _T_4803_re;
    _T_4804_im <= _T_4803_im;
    _T_4805_re <= _T_4804_re;
    _T_4805_im <= _T_4804_im;
    _T_4811_re <= Switch_1_io_out1_re;
    _T_4811_im <= Switch_1_io_out1_im;
    _T_4812_re <= _T_4811_re;
    _T_4812_im <= _T_4811_im;
    _T_4813_re <= _T_4812_re;
    _T_4813_im <= _T_4812_im;
    _T_4814_re <= _T_4813_re;
    _T_4814_im <= _T_4813_im;
    _T_4815_re <= _T_4814_re;
    _T_4815_im <= _T_4814_im;
    _T_4816_re <= _T_4815_re;
    _T_4816_im <= _T_4815_im;
    _T_4817_re <= _T_4816_re;
    _T_4817_im <= _T_4816_im;
    _T_4818_re <= _T_4817_re;
    _T_4818_im <= _T_4817_im;
    _T_4819_re <= _T_4818_re;
    _T_4819_im <= _T_4818_im;
    _T_4820_re <= _T_4819_re;
    _T_4820_im <= _T_4819_im;
    _T_4821_re <= _T_4820_re;
    _T_4821_im <= _T_4820_im;
    _T_4822_re <= _T_4821_re;
    _T_4822_im <= _T_4821_im;
    _T_4823_re <= _T_4822_re;
    _T_4823_im <= _T_4822_im;
    _T_4824_re <= _T_4823_re;
    _T_4824_im <= _T_4823_im;
    _T_4825_re <= _T_4824_re;
    _T_4825_im <= _T_4824_im;
    _T_4826_re <= _T_4825_re;
    _T_4826_im <= _T_4825_im;
    _T_4827_re <= _T_4826_re;
    _T_4827_im <= _T_4826_im;
    _T_4828_re <= _T_4827_re;
    _T_4828_im <= _T_4827_im;
    _T_4829_re <= _T_4828_re;
    _T_4829_im <= _T_4828_im;
    _T_4830_re <= _T_4829_re;
    _T_4830_im <= _T_4829_im;
    _T_4831_re <= _T_4830_re;
    _T_4831_im <= _T_4830_im;
    _T_4832_re <= _T_4831_re;
    _T_4832_im <= _T_4831_im;
    _T_4833_re <= _T_4832_re;
    _T_4833_im <= _T_4832_im;
    _T_4834_re <= _T_4833_re;
    _T_4834_im <= _T_4833_im;
    _T_4835_re <= _T_4834_re;
    _T_4835_im <= _T_4834_im;
    _T_4836_re <= _T_4835_re;
    _T_4836_im <= _T_4835_im;
    _T_4837_re <= _T_4836_re;
    _T_4837_im <= _T_4836_im;
    _T_4838_re <= _T_4837_re;
    _T_4838_im <= _T_4837_im;
    _T_4839_re <= _T_4838_re;
    _T_4839_im <= _T_4838_im;
    _T_4840_re <= _T_4839_re;
    _T_4840_im <= _T_4839_im;
    _T_4841_re <= _T_4840_re;
    _T_4841_im <= _T_4840_im;
    _T_4842_re <= _T_4841_re;
    _T_4842_im <= _T_4841_im;
    _T_4843_re <= _T_4842_re;
    _T_4843_im <= _T_4842_im;
    _T_4844_re <= _T_4843_re;
    _T_4844_im <= _T_4843_im;
    _T_4845_re <= _T_4844_re;
    _T_4845_im <= _T_4844_im;
    _T_4846_re <= _T_4845_re;
    _T_4846_im <= _T_4845_im;
    _T_4847_re <= _T_4846_re;
    _T_4847_im <= _T_4846_im;
    _T_4848_re <= _T_4847_re;
    _T_4848_im <= _T_4847_im;
    _T_4849_re <= _T_4848_re;
    _T_4849_im <= _T_4848_im;
    _T_4850_re <= _T_4849_re;
    _T_4850_im <= _T_4849_im;
    _T_4851_re <= _T_4850_re;
    _T_4851_im <= _T_4850_im;
    _T_4852_re <= _T_4851_re;
    _T_4852_im <= _T_4851_im;
    _T_4853_re <= _T_4852_re;
    _T_4853_im <= _T_4852_im;
    _T_4854_re <= _T_4853_re;
    _T_4854_im <= _T_4853_im;
    _T_4855_re <= _T_4854_re;
    _T_4855_im <= _T_4854_im;
    _T_4856_re <= _T_4855_re;
    _T_4856_im <= _T_4855_im;
    _T_4857_re <= _T_4856_re;
    _T_4857_im <= _T_4856_im;
    _T_4858_re <= _T_4857_re;
    _T_4858_im <= _T_4857_im;
    _T_4859_re <= _T_4858_re;
    _T_4859_im <= _T_4858_im;
    _T_4860_re <= _T_4859_re;
    _T_4860_im <= _T_4859_im;
    _T_4861_re <= _T_4860_re;
    _T_4861_im <= _T_4860_im;
    _T_4862_re <= _T_4861_re;
    _T_4862_im <= _T_4861_im;
    _T_4863_re <= _T_4862_re;
    _T_4863_im <= _T_4862_im;
    _T_4864_re <= _T_4863_re;
    _T_4864_im <= _T_4863_im;
    _T_4865_re <= _T_4864_re;
    _T_4865_im <= _T_4864_im;
    _T_4866_re <= _T_4865_re;
    _T_4866_im <= _T_4865_im;
    _T_4867_re <= _T_4866_re;
    _T_4867_im <= _T_4866_im;
    _T_4868_re <= _T_4867_re;
    _T_4868_im <= _T_4867_im;
    _T_4869_re <= _T_4868_re;
    _T_4869_im <= _T_4868_im;
    _T_4870_re <= _T_4869_re;
    _T_4870_im <= _T_4869_im;
    _T_4871_re <= _T_4870_re;
    _T_4871_im <= _T_4870_im;
    _T_4872_re <= _T_4871_re;
    _T_4872_im <= _T_4871_im;
    _T_4873_re <= _T_4872_re;
    _T_4873_im <= _T_4872_im;
    _T_4874_re <= _T_4873_re;
    _T_4874_im <= _T_4873_im;
    _T_4875_re <= _T_4874_re;
    _T_4875_im <= _T_4874_im;
    _T_4876_re <= _T_4875_re;
    _T_4876_im <= _T_4875_im;
    _T_4877_re <= _T_4876_re;
    _T_4877_im <= _T_4876_im;
    _T_4878_re <= _T_4877_re;
    _T_4878_im <= _T_4877_im;
    _T_4879_re <= _T_4878_re;
    _T_4879_im <= _T_4878_im;
    _T_4880_re <= _T_4879_re;
    _T_4880_im <= _T_4879_im;
    _T_4881_re <= _T_4880_re;
    _T_4881_im <= _T_4880_im;
    _T_4882_re <= _T_4881_re;
    _T_4882_im <= _T_4881_im;
    _T_4883_re <= _T_4882_re;
    _T_4883_im <= _T_4882_im;
    _T_4884_re <= _T_4883_re;
    _T_4884_im <= _T_4883_im;
    _T_4885_re <= _T_4884_re;
    _T_4885_im <= _T_4884_im;
    _T_4886_re <= _T_4885_re;
    _T_4886_im <= _T_4885_im;
    _T_4887_re <= _T_4886_re;
    _T_4887_im <= _T_4886_im;
    _T_4888_re <= _T_4887_re;
    _T_4888_im <= _T_4887_im;
    _T_4889_re <= _T_4888_re;
    _T_4889_im <= _T_4888_im;
    _T_4890_re <= _T_4889_re;
    _T_4890_im <= _T_4889_im;
    _T_4891_re <= _T_4890_re;
    _T_4891_im <= _T_4890_im;
    _T_4892_re <= _T_4891_re;
    _T_4892_im <= _T_4891_im;
    _T_4893_re <= _T_4892_re;
    _T_4893_im <= _T_4892_im;
    _T_4894_re <= _T_4893_re;
    _T_4894_im <= _T_4893_im;
    _T_4895_re <= _T_4894_re;
    _T_4895_im <= _T_4894_im;
    _T_4896_re <= _T_4895_re;
    _T_4896_im <= _T_4895_im;
    _T_4897_re <= _T_4896_re;
    _T_4897_im <= _T_4896_im;
    _T_4898_re <= _T_4897_re;
    _T_4898_im <= _T_4897_im;
    _T_4899_re <= _T_4898_re;
    _T_4899_im <= _T_4898_im;
    _T_4900_re <= _T_4899_re;
    _T_4900_im <= _T_4899_im;
    _T_4901_re <= _T_4900_re;
    _T_4901_im <= _T_4900_im;
    _T_4902_re <= _T_4901_re;
    _T_4902_im <= _T_4901_im;
    _T_4903_re <= _T_4902_re;
    _T_4903_im <= _T_4902_im;
    _T_4904_re <= _T_4903_re;
    _T_4904_im <= _T_4903_im;
    _T_4905_re <= _T_4904_re;
    _T_4905_im <= _T_4904_im;
    _T_4906_re <= _T_4905_re;
    _T_4906_im <= _T_4905_im;
    _T_4907_re <= _T_4906_re;
    _T_4907_im <= _T_4906_im;
    _T_4908_re <= _T_4907_re;
    _T_4908_im <= _T_4907_im;
    _T_4909_re <= _T_4908_re;
    _T_4909_im <= _T_4908_im;
    _T_4910_re <= _T_4909_re;
    _T_4910_im <= _T_4909_im;
    _T_4911_re <= _T_4910_re;
    _T_4911_im <= _T_4910_im;
    _T_4912_re <= _T_4911_re;
    _T_4912_im <= _T_4911_im;
    _T_4913_re <= _T_4912_re;
    _T_4913_im <= _T_4912_im;
    _T_4914_re <= _T_4913_re;
    _T_4914_im <= _T_4913_im;
    _T_4915_re <= _T_4914_re;
    _T_4915_im <= _T_4914_im;
    _T_4916_re <= _T_4915_re;
    _T_4916_im <= _T_4915_im;
    _T_4917_re <= _T_4916_re;
    _T_4917_im <= _T_4916_im;
    _T_4918_re <= _T_4917_re;
    _T_4918_im <= _T_4917_im;
    _T_4919_re <= _T_4918_re;
    _T_4919_im <= _T_4918_im;
    _T_4920_re <= _T_4919_re;
    _T_4920_im <= _T_4919_im;
    _T_4921_re <= _T_4920_re;
    _T_4921_im <= _T_4920_im;
    _T_4922_re <= _T_4921_re;
    _T_4922_im <= _T_4921_im;
    _T_4923_re <= _T_4922_re;
    _T_4923_im <= _T_4922_im;
    _T_4924_re <= _T_4923_re;
    _T_4924_im <= _T_4923_im;
    _T_4925_re <= _T_4924_re;
    _T_4925_im <= _T_4924_im;
    _T_4926_re <= _T_4925_re;
    _T_4926_im <= _T_4925_im;
    _T_4927_re <= _T_4926_re;
    _T_4927_im <= _T_4926_im;
    _T_4928_re <= _T_4927_re;
    _T_4928_im <= _T_4927_im;
    _T_4929_re <= _T_4928_re;
    _T_4929_im <= _T_4928_im;
    _T_4930_re <= _T_4929_re;
    _T_4930_im <= _T_4929_im;
    _T_4931_re <= _T_4930_re;
    _T_4931_im <= _T_4930_im;
    _T_4932_re <= _T_4931_re;
    _T_4932_im <= _T_4931_im;
    _T_4933_re <= _T_4932_re;
    _T_4933_im <= _T_4932_im;
    _T_4934_re <= _T_4933_re;
    _T_4934_im <= _T_4933_im;
    _T_4935_re <= _T_4934_re;
    _T_4935_im <= _T_4934_im;
    _T_4936_re <= _T_4935_re;
    _T_4936_im <= _T_4935_im;
    _T_4937_re <= _T_4936_re;
    _T_4937_im <= _T_4936_im;
    _T_4938_re <= _T_4937_re;
    _T_4938_im <= _T_4937_im;
    _T_4939_re <= _T_4938_re;
    _T_4939_im <= _T_4938_im;
    _T_4940_re <= _T_4939_re;
    _T_4940_im <= _T_4939_im;
    _T_4941_re <= _T_4940_re;
    _T_4941_im <= _T_4940_im;
    _T_4942_re <= _T_4941_re;
    _T_4942_im <= _T_4941_im;
    _T_4943_re <= _T_4942_re;
    _T_4943_im <= _T_4942_im;
    _T_4944_re <= _T_4943_re;
    _T_4944_im <= _T_4943_im;
    _T_4945_re <= _T_4944_re;
    _T_4945_im <= _T_4944_im;
    _T_4946_re <= _T_4945_re;
    _T_4946_im <= _T_4945_im;
    _T_4947_re <= _T_4946_re;
    _T_4947_im <= _T_4946_im;
    _T_4948_re <= _T_4947_re;
    _T_4948_im <= _T_4947_im;
    _T_4949_re <= _T_4948_re;
    _T_4949_im <= _T_4948_im;
    _T_4950_re <= _T_4949_re;
    _T_4950_im <= _T_4949_im;
    _T_4951_re <= _T_4950_re;
    _T_4951_im <= _T_4950_im;
    _T_4952_re <= _T_4951_re;
    _T_4952_im <= _T_4951_im;
    _T_4953_re <= _T_4952_re;
    _T_4953_im <= _T_4952_im;
    _T_4954_re <= _T_4953_re;
    _T_4954_im <= _T_4953_im;
    _T_4955_re <= _T_4954_re;
    _T_4955_im <= _T_4954_im;
    _T_4956_re <= _T_4955_re;
    _T_4956_im <= _T_4955_im;
    _T_4957_re <= _T_4956_re;
    _T_4957_im <= _T_4956_im;
    _T_4958_re <= _T_4957_re;
    _T_4958_im <= _T_4957_im;
    _T_4959_re <= _T_4958_re;
    _T_4959_im <= _T_4958_im;
    _T_4960_re <= _T_4959_re;
    _T_4960_im <= _T_4959_im;
    _T_4961_re <= _T_4960_re;
    _T_4961_im <= _T_4960_im;
    _T_4962_re <= _T_4961_re;
    _T_4962_im <= _T_4961_im;
    _T_4963_re <= _T_4962_re;
    _T_4963_im <= _T_4962_im;
    _T_4964_re <= _T_4963_re;
    _T_4964_im <= _T_4963_im;
    _T_4965_re <= _T_4964_re;
    _T_4965_im <= _T_4964_im;
    _T_4966_re <= _T_4965_re;
    _T_4966_im <= _T_4965_im;
    _T_4967_re <= _T_4966_re;
    _T_4967_im <= _T_4966_im;
    _T_4968_re <= _T_4967_re;
    _T_4968_im <= _T_4967_im;
    _T_4969_re <= _T_4968_re;
    _T_4969_im <= _T_4968_im;
    _T_4970_re <= _T_4969_re;
    _T_4970_im <= _T_4969_im;
    _T_4971_re <= _T_4970_re;
    _T_4971_im <= _T_4970_im;
    _T_4972_re <= _T_4971_re;
    _T_4972_im <= _T_4971_im;
    _T_4973_re <= _T_4972_re;
    _T_4973_im <= _T_4972_im;
    _T_4974_re <= _T_4973_re;
    _T_4974_im <= _T_4973_im;
    _T_4975_re <= _T_4974_re;
    _T_4975_im <= _T_4974_im;
    _T_4976_re <= _T_4975_re;
    _T_4976_im <= _T_4975_im;
    _T_4977_re <= _T_4976_re;
    _T_4977_im <= _T_4976_im;
    _T_4978_re <= _T_4977_re;
    _T_4978_im <= _T_4977_im;
    _T_4979_re <= _T_4978_re;
    _T_4979_im <= _T_4978_im;
    _T_4980_re <= _T_4979_re;
    _T_4980_im <= _T_4979_im;
    _T_4981_re <= _T_4980_re;
    _T_4981_im <= _T_4980_im;
    _T_4982_re <= _T_4981_re;
    _T_4982_im <= _T_4981_im;
    _T_4983_re <= _T_4982_re;
    _T_4983_im <= _T_4982_im;
    _T_4984_re <= _T_4983_re;
    _T_4984_im <= _T_4983_im;
    _T_4985_re <= _T_4984_re;
    _T_4985_im <= _T_4984_im;
    _T_4986_re <= _T_4985_re;
    _T_4986_im <= _T_4985_im;
    _T_4987_re <= _T_4986_re;
    _T_4987_im <= _T_4986_im;
    _T_4988_re <= _T_4987_re;
    _T_4988_im <= _T_4987_im;
    _T_4989_re <= _T_4988_re;
    _T_4989_im <= _T_4988_im;
    _T_4990_re <= _T_4989_re;
    _T_4990_im <= _T_4989_im;
    _T_4991_re <= _T_4990_re;
    _T_4991_im <= _T_4990_im;
    _T_4992_re <= _T_4991_re;
    _T_4992_im <= _T_4991_im;
    _T_4993_re <= _T_4992_re;
    _T_4993_im <= _T_4992_im;
    _T_4994_re <= _T_4993_re;
    _T_4994_im <= _T_4993_im;
    _T_4995_re <= _T_4994_re;
    _T_4995_im <= _T_4994_im;
    _T_4996_re <= _T_4995_re;
    _T_4996_im <= _T_4995_im;
    _T_4997_re <= _T_4996_re;
    _T_4997_im <= _T_4996_im;
    _T_4998_re <= _T_4997_re;
    _T_4998_im <= _T_4997_im;
    _T_4999_re <= _T_4998_re;
    _T_4999_im <= _T_4998_im;
    _T_5000_re <= _T_4999_re;
    _T_5000_im <= _T_4999_im;
    _T_5001_re <= _T_5000_re;
    _T_5001_im <= _T_5000_im;
    _T_5002_re <= _T_5001_re;
    _T_5002_im <= _T_5001_im;
    _T_5003_re <= _T_5002_re;
    _T_5003_im <= _T_5002_im;
    _T_5004_re <= _T_5003_re;
    _T_5004_im <= _T_5003_im;
    _T_5005_re <= _T_5004_re;
    _T_5005_im <= _T_5004_im;
    _T_5006_re <= _T_5005_re;
    _T_5006_im <= _T_5005_im;
    _T_5007_re <= _T_5006_re;
    _T_5007_im <= _T_5006_im;
    _T_5008_re <= _T_5007_re;
    _T_5008_im <= _T_5007_im;
    _T_5009_re <= _T_5008_re;
    _T_5009_im <= _T_5008_im;
    _T_5010_re <= _T_5009_re;
    _T_5010_im <= _T_5009_im;
    _T_5011_re <= _T_5010_re;
    _T_5011_im <= _T_5010_im;
    _T_5012_re <= _T_5011_re;
    _T_5012_im <= _T_5011_im;
    _T_5013_re <= _T_5012_re;
    _T_5013_im <= _T_5012_im;
    _T_5014_re <= _T_5013_re;
    _T_5014_im <= _T_5013_im;
    _T_5015_re <= _T_5014_re;
    _T_5015_im <= _T_5014_im;
    _T_5016_re <= _T_5015_re;
    _T_5016_im <= _T_5015_im;
    _T_5017_re <= _T_5016_re;
    _T_5017_im <= _T_5016_im;
    _T_5018_re <= _T_5017_re;
    _T_5018_im <= _T_5017_im;
    _T_5019_re <= _T_5018_re;
    _T_5019_im <= _T_5018_im;
    _T_5020_re <= _T_5019_re;
    _T_5020_im <= _T_5019_im;
    _T_5021_re <= _T_5020_re;
    _T_5021_im <= _T_5020_im;
    _T_5022_re <= _T_5021_re;
    _T_5022_im <= _T_5021_im;
    _T_5023_re <= _T_5022_re;
    _T_5023_im <= _T_5022_im;
    _T_5024_re <= _T_5023_re;
    _T_5024_im <= _T_5023_im;
    _T_5025_re <= _T_5024_re;
    _T_5025_im <= _T_5024_im;
    _T_5026_re <= _T_5025_re;
    _T_5026_im <= _T_5025_im;
    _T_5027_re <= _T_5026_re;
    _T_5027_im <= _T_5026_im;
    _T_5028_re <= _T_5027_re;
    _T_5028_im <= _T_5027_im;
    _T_5029_re <= _T_5028_re;
    _T_5029_im <= _T_5028_im;
    _T_5030_re <= _T_5029_re;
    _T_5030_im <= _T_5029_im;
    _T_5031_re <= _T_5030_re;
    _T_5031_im <= _T_5030_im;
    _T_5032_re <= _T_5031_re;
    _T_5032_im <= _T_5031_im;
    _T_5033_re <= _T_5032_re;
    _T_5033_im <= _T_5032_im;
    _T_5034_re <= _T_5033_re;
    _T_5034_im <= _T_5033_im;
    _T_5035_re <= _T_5034_re;
    _T_5035_im <= _T_5034_im;
    _T_5036_re <= _T_5035_re;
    _T_5036_im <= _T_5035_im;
    _T_5037_re <= _T_5036_re;
    _T_5037_im <= _T_5036_im;
    _T_5038_re <= _T_5037_re;
    _T_5038_im <= _T_5037_im;
    _T_5039_re <= _T_5038_re;
    _T_5039_im <= _T_5038_im;
    _T_5040_re <= _T_5039_re;
    _T_5040_im <= _T_5039_im;
    _T_5041_re <= _T_5040_re;
    _T_5041_im <= _T_5040_im;
    _T_5042_re <= _T_5041_re;
    _T_5042_im <= _T_5041_im;
    _T_5043_re <= _T_5042_re;
    _T_5043_im <= _T_5042_im;
    _T_5044_re <= _T_5043_re;
    _T_5044_im <= _T_5043_im;
    _T_5045_re <= _T_5044_re;
    _T_5045_im <= _T_5044_im;
    _T_5046_re <= _T_5045_re;
    _T_5046_im <= _T_5045_im;
    _T_5047_re <= _T_5046_re;
    _T_5047_im <= _T_5046_im;
    _T_5048_re <= _T_5047_re;
    _T_5048_im <= _T_5047_im;
    _T_5049_re <= _T_5048_re;
    _T_5049_im <= _T_5048_im;
    _T_5050_re <= _T_5049_re;
    _T_5050_im <= _T_5049_im;
    _T_5051_re <= _T_5050_re;
    _T_5051_im <= _T_5050_im;
    _T_5052_re <= _T_5051_re;
    _T_5052_im <= _T_5051_im;
    _T_5053_re <= _T_5052_re;
    _T_5053_im <= _T_5052_im;
    _T_5054_re <= _T_5053_re;
    _T_5054_im <= _T_5053_im;
    _T_5055_re <= _T_5054_re;
    _T_5055_im <= _T_5054_im;
    _T_5056_re <= _T_5055_re;
    _T_5056_im <= _T_5055_im;
    _T_5057_re <= _T_5056_re;
    _T_5057_im <= _T_5056_im;
    _T_5058_re <= _T_5057_re;
    _T_5058_im <= _T_5057_im;
    _T_5059_re <= _T_5058_re;
    _T_5059_im <= _T_5058_im;
    _T_5060_re <= _T_5059_re;
    _T_5060_im <= _T_5059_im;
    _T_5061_re <= _T_5060_re;
    _T_5061_im <= _T_5060_im;
    _T_5062_re <= _T_5061_re;
    _T_5062_im <= _T_5061_im;
    _T_5063_re <= _T_5062_re;
    _T_5063_im <= _T_5062_im;
    _T_5064_re <= _T_5063_re;
    _T_5064_im <= _T_5063_im;
    _T_5065_re <= _T_5064_re;
    _T_5065_im <= _T_5064_im;
    _T_5066_re <= _T_5065_re;
    _T_5066_im <= _T_5065_im;
    _T_5067_re <= _T_5066_re;
    _T_5067_im <= _T_5066_im;
    _T_5068_re <= _T_5067_re;
    _T_5068_im <= _T_5067_im;
    _T_5069_re <= _T_5068_re;
    _T_5069_im <= _T_5068_im;
    _T_5070_re <= _T_5069_re;
    _T_5070_im <= _T_5069_im;
    _T_5071_re <= _T_5070_re;
    _T_5071_im <= _T_5070_im;
    _T_5072_re <= _T_5071_re;
    _T_5072_im <= _T_5071_im;
    _T_5073_re <= _T_5072_re;
    _T_5073_im <= _T_5072_im;
    _T_5074_re <= _T_5073_re;
    _T_5074_im <= _T_5073_im;
    _T_5075_re <= _T_5074_re;
    _T_5075_im <= _T_5074_im;
    _T_5076_re <= _T_5075_re;
    _T_5076_im <= _T_5075_im;
    _T_5077_re <= _T_5076_re;
    _T_5077_im <= _T_5076_im;
    _T_5078_re <= _T_5077_re;
    _T_5078_im <= _T_5077_im;
    _T_5079_re <= _T_5078_re;
    _T_5079_im <= _T_5078_im;
    _T_5080_re <= _T_5079_re;
    _T_5080_im <= _T_5079_im;
    _T_5081_re <= _T_5080_re;
    _T_5081_im <= _T_5080_im;
    _T_5082_re <= _T_5081_re;
    _T_5082_im <= _T_5081_im;
    _T_5083_re <= _T_5082_re;
    _T_5083_im <= _T_5082_im;
    _T_5084_re <= _T_5083_re;
    _T_5084_im <= _T_5083_im;
    _T_5085_re <= _T_5084_re;
    _T_5085_im <= _T_5084_im;
    _T_5086_re <= _T_5085_re;
    _T_5086_im <= _T_5085_im;
    _T_5087_re <= _T_5086_re;
    _T_5087_im <= _T_5086_im;
    _T_5088_re <= _T_5087_re;
    _T_5088_im <= _T_5087_im;
    _T_5089_re <= _T_5088_re;
    _T_5089_im <= _T_5088_im;
    _T_5090_re <= _T_5089_re;
    _T_5090_im <= _T_5089_im;
    _T_5091_re <= _T_5090_re;
    _T_5091_im <= _T_5090_im;
    _T_5092_re <= _T_5091_re;
    _T_5092_im <= _T_5091_im;
    _T_5093_re <= _T_5092_re;
    _T_5093_im <= _T_5092_im;
    _T_5094_re <= _T_5093_re;
    _T_5094_im <= _T_5093_im;
    _T_5095_re <= _T_5094_re;
    _T_5095_im <= _T_5094_im;
    _T_5096_re <= _T_5095_re;
    _T_5096_im <= _T_5095_im;
    _T_5097_re <= _T_5096_re;
    _T_5097_im <= _T_5096_im;
    _T_5098_re <= _T_5097_re;
    _T_5098_im <= _T_5097_im;
    _T_5099_re <= _T_5098_re;
    _T_5099_im <= _T_5098_im;
    _T_5100_re <= _T_5099_re;
    _T_5100_im <= _T_5099_im;
    _T_5101_re <= _T_5100_re;
    _T_5101_im <= _T_5100_im;
    _T_5102_re <= _T_5101_re;
    _T_5102_im <= _T_5101_im;
    _T_5103_re <= _T_5102_re;
    _T_5103_im <= _T_5102_im;
    _T_5104_re <= _T_5103_re;
    _T_5104_im <= _T_5103_im;
    _T_5105_re <= _T_5104_re;
    _T_5105_im <= _T_5104_im;
    _T_5106_re <= _T_5105_re;
    _T_5106_im <= _T_5105_im;
    _T_5107_re <= _T_5106_re;
    _T_5107_im <= _T_5106_im;
    _T_5108_re <= _T_5107_re;
    _T_5108_im <= _T_5107_im;
    _T_5109_re <= _T_5108_re;
    _T_5109_im <= _T_5108_im;
    _T_5110_re <= _T_5109_re;
    _T_5110_im <= _T_5109_im;
    _T_5111_re <= _T_5110_re;
    _T_5111_im <= _T_5110_im;
    _T_5112_re <= _T_5111_re;
    _T_5112_im <= _T_5111_im;
    _T_5113_re <= _T_5112_re;
    _T_5113_im <= _T_5112_im;
    _T_5114_re <= _T_5113_re;
    _T_5114_im <= _T_5113_im;
    _T_5115_re <= _T_5114_re;
    _T_5115_im <= _T_5114_im;
    _T_5116_re <= _T_5115_re;
    _T_5116_im <= _T_5115_im;
    _T_5117_re <= _T_5116_re;
    _T_5117_im <= _T_5116_im;
    _T_5118_re <= _T_5117_re;
    _T_5118_im <= _T_5117_im;
    _T_5119_re <= _T_5118_re;
    _T_5119_im <= _T_5118_im;
    _T_5120_re <= _T_5119_re;
    _T_5120_im <= _T_5119_im;
    _T_5121_re <= _T_5120_re;
    _T_5121_im <= _T_5120_im;
    _T_5122_re <= _T_5121_re;
    _T_5122_im <= _T_5121_im;
    _T_5123_re <= _T_5122_re;
    _T_5123_im <= _T_5122_im;
    _T_5124_re <= _T_5123_re;
    _T_5124_im <= _T_5123_im;
    _T_5125_re <= _T_5124_re;
    _T_5125_im <= _T_5124_im;
    _T_5126_re <= _T_5125_re;
    _T_5126_im <= _T_5125_im;
    _T_5127_re <= _T_5126_re;
    _T_5127_im <= _T_5126_im;
    _T_5128_re <= _T_5127_re;
    _T_5128_im <= _T_5127_im;
    _T_5129_re <= _T_5128_re;
    _T_5129_im <= _T_5128_im;
    _T_5130_re <= _T_5129_re;
    _T_5130_im <= _T_5129_im;
    _T_5131_re <= _T_5130_re;
    _T_5131_im <= _T_5130_im;
    _T_5132_re <= _T_5131_re;
    _T_5132_im <= _T_5131_im;
    _T_5133_re <= _T_5132_re;
    _T_5133_im <= _T_5132_im;
    _T_5134_re <= _T_5133_re;
    _T_5134_im <= _T_5133_im;
    _T_5135_re <= _T_5134_re;
    _T_5135_im <= _T_5134_im;
    _T_5136_re <= _T_5135_re;
    _T_5136_im <= _T_5135_im;
    _T_5137_re <= _T_5136_re;
    _T_5137_im <= _T_5136_im;
    _T_5138_re <= _T_5137_re;
    _T_5138_im <= _T_5137_im;
    _T_5139_re <= _T_5138_re;
    _T_5139_im <= _T_5138_im;
    _T_5140_re <= _T_5139_re;
    _T_5140_im <= _T_5139_im;
    _T_5141_re <= _T_5140_re;
    _T_5141_im <= _T_5140_im;
    _T_5142_re <= _T_5141_re;
    _T_5142_im <= _T_5141_im;
    _T_5143_re <= _T_5142_re;
    _T_5143_im <= _T_5142_im;
    _T_5144_re <= _T_5143_re;
    _T_5144_im <= _T_5143_im;
    _T_5145_re <= _T_5144_re;
    _T_5145_im <= _T_5144_im;
    _T_5146_re <= _T_5145_re;
    _T_5146_im <= _T_5145_im;
    _T_5147_re <= _T_5146_re;
    _T_5147_im <= _T_5146_im;
    _T_5148_re <= _T_5147_re;
    _T_5148_im <= _T_5147_im;
    _T_5149_re <= _T_5148_re;
    _T_5149_im <= _T_5148_im;
    _T_5150_re <= _T_5149_re;
    _T_5150_im <= _T_5149_im;
    _T_5151_re <= _T_5150_re;
    _T_5151_im <= _T_5150_im;
    _T_5152_re <= _T_5151_re;
    _T_5152_im <= _T_5151_im;
    _T_5153_re <= _T_5152_re;
    _T_5153_im <= _T_5152_im;
    _T_5154_re <= _T_5153_re;
    _T_5154_im <= _T_5153_im;
    _T_5155_re <= _T_5154_re;
    _T_5155_im <= _T_5154_im;
    _T_5156_re <= _T_5155_re;
    _T_5156_im <= _T_5155_im;
    _T_5157_re <= _T_5156_re;
    _T_5157_im <= _T_5156_im;
    _T_5158_re <= _T_5157_re;
    _T_5158_im <= _T_5157_im;
    _T_5159_re <= _T_5158_re;
    _T_5159_im <= _T_5158_im;
    _T_5160_re <= _T_5159_re;
    _T_5160_im <= _T_5159_im;
    _T_5161_re <= _T_5160_re;
    _T_5161_im <= _T_5160_im;
    _T_5162_re <= _T_5161_re;
    _T_5162_im <= _T_5161_im;
    _T_5163_re <= _T_5162_re;
    _T_5163_im <= _T_5162_im;
    _T_5164_re <= _T_5163_re;
    _T_5164_im <= _T_5163_im;
    _T_5165_re <= _T_5164_re;
    _T_5165_im <= _T_5164_im;
    _T_5166_re <= _T_5165_re;
    _T_5166_im <= _T_5165_im;
    _T_5167_re <= _T_5166_re;
    _T_5167_im <= _T_5166_im;
    _T_5168_re <= _T_5167_re;
    _T_5168_im <= _T_5167_im;
    _T_5169_re <= _T_5168_re;
    _T_5169_im <= _T_5168_im;
    _T_5170_re <= _T_5169_re;
    _T_5170_im <= _T_5169_im;
    _T_5171_re <= _T_5170_re;
    _T_5171_im <= _T_5170_im;
    _T_5172_re <= _T_5171_re;
    _T_5172_im <= _T_5171_im;
    _T_5173_re <= _T_5172_re;
    _T_5173_im <= _T_5172_im;
    _T_5174_re <= _T_5173_re;
    _T_5174_im <= _T_5173_im;
    _T_5175_re <= _T_5174_re;
    _T_5175_im <= _T_5174_im;
    _T_5176_re <= _T_5175_re;
    _T_5176_im <= _T_5175_im;
    _T_5177_re <= _T_5176_re;
    _T_5177_im <= _T_5176_im;
    _T_5178_re <= _T_5177_re;
    _T_5178_im <= _T_5177_im;
    _T_5179_re <= _T_5178_re;
    _T_5179_im <= _T_5178_im;
    _T_5180_re <= _T_5179_re;
    _T_5180_im <= _T_5179_im;
    _T_5181_re <= _T_5180_re;
    _T_5181_im <= _T_5180_im;
    _T_5182_re <= _T_5181_re;
    _T_5182_im <= _T_5181_im;
    _T_5183_re <= _T_5182_re;
    _T_5183_im <= _T_5182_im;
    _T_5184_re <= _T_5183_re;
    _T_5184_im <= _T_5183_im;
    _T_5185_re <= _T_5184_re;
    _T_5185_im <= _T_5184_im;
    _T_5186_re <= _T_5185_re;
    _T_5186_im <= _T_5185_im;
    _T_5187_re <= _T_5186_re;
    _T_5187_im <= _T_5186_im;
    _T_5188_re <= _T_5187_re;
    _T_5188_im <= _T_5187_im;
    _T_5189_re <= _T_5188_re;
    _T_5189_im <= _T_5188_im;
    _T_5190_re <= _T_5189_re;
    _T_5190_im <= _T_5189_im;
    _T_5191_re <= _T_5190_re;
    _T_5191_im <= _T_5190_im;
    _T_5192_re <= _T_5191_re;
    _T_5192_im <= _T_5191_im;
    _T_5193_re <= _T_5192_re;
    _T_5193_im <= _T_5192_im;
    _T_5194_re <= _T_5193_re;
    _T_5194_im <= _T_5193_im;
    _T_5195_re <= _T_5194_re;
    _T_5195_im <= _T_5194_im;
    _T_5196_re <= _T_5195_re;
    _T_5196_im <= _T_5195_im;
    _T_5197_re <= _T_5196_re;
    _T_5197_im <= _T_5196_im;
    _T_5198_re <= _T_5197_re;
    _T_5198_im <= _T_5197_im;
    _T_5199_re <= _T_5198_re;
    _T_5199_im <= _T_5198_im;
    _T_5200_re <= _T_5199_re;
    _T_5200_im <= _T_5199_im;
    _T_5201_re <= _T_5200_re;
    _T_5201_im <= _T_5200_im;
    _T_5202_re <= _T_5201_re;
    _T_5202_im <= _T_5201_im;
    _T_5203_re <= _T_5202_re;
    _T_5203_im <= _T_5202_im;
    _T_5204_re <= _T_5203_re;
    _T_5204_im <= _T_5203_im;
    _T_5205_re <= _T_5204_re;
    _T_5205_im <= _T_5204_im;
    _T_5206_re <= _T_5205_re;
    _T_5206_im <= _T_5205_im;
    _T_5207_re <= _T_5206_re;
    _T_5207_im <= _T_5206_im;
    _T_5208_re <= _T_5207_re;
    _T_5208_im <= _T_5207_im;
    _T_5209_re <= _T_5208_re;
    _T_5209_im <= _T_5208_im;
    _T_5210_re <= _T_5209_re;
    _T_5210_im <= _T_5209_im;
    _T_5211_re <= _T_5210_re;
    _T_5211_im <= _T_5210_im;
    _T_5212_re <= _T_5211_re;
    _T_5212_im <= _T_5211_im;
    _T_5213_re <= _T_5212_re;
    _T_5213_im <= _T_5212_im;
    _T_5214_re <= _T_5213_re;
    _T_5214_im <= _T_5213_im;
    _T_5215_re <= _T_5214_re;
    _T_5215_im <= _T_5214_im;
    _T_5216_re <= _T_5215_re;
    _T_5216_im <= _T_5215_im;
    _T_5217_re <= _T_5216_re;
    _T_5217_im <= _T_5216_im;
    _T_5218_re <= _T_5217_re;
    _T_5218_im <= _T_5217_im;
    _T_5219_re <= _T_5218_re;
    _T_5219_im <= _T_5218_im;
    _T_5220_re <= _T_5219_re;
    _T_5220_im <= _T_5219_im;
    _T_5221_re <= _T_5220_re;
    _T_5221_im <= _T_5220_im;
    _T_5222_re <= _T_5221_re;
    _T_5222_im <= _T_5221_im;
    _T_5223_re <= _T_5222_re;
    _T_5223_im <= _T_5222_im;
    _T_5224_re <= _T_5223_re;
    _T_5224_im <= _T_5223_im;
    _T_5225_re <= _T_5224_re;
    _T_5225_im <= _T_5224_im;
    _T_5226_re <= _T_5225_re;
    _T_5226_im <= _T_5225_im;
    _T_5227_re <= _T_5226_re;
    _T_5227_im <= _T_5226_im;
    _T_5228_re <= _T_5227_re;
    _T_5228_im <= _T_5227_im;
    _T_5229_re <= _T_5228_re;
    _T_5229_im <= _T_5228_im;
    _T_5230_re <= _T_5229_re;
    _T_5230_im <= _T_5229_im;
    _T_5231_re <= _T_5230_re;
    _T_5231_im <= _T_5230_im;
    _T_5232_re <= _T_5231_re;
    _T_5232_im <= _T_5231_im;
    _T_5233_re <= _T_5232_re;
    _T_5233_im <= _T_5232_im;
    _T_5234_re <= _T_5233_re;
    _T_5234_im <= _T_5233_im;
    _T_5235_re <= _T_5234_re;
    _T_5235_im <= _T_5234_im;
    _T_5236_re <= _T_5235_re;
    _T_5236_im <= _T_5235_im;
    _T_5237_re <= _T_5236_re;
    _T_5237_im <= _T_5236_im;
    _T_5238_re <= _T_5237_re;
    _T_5238_im <= _T_5237_im;
    _T_5239_re <= _T_5238_re;
    _T_5239_im <= _T_5238_im;
    _T_5240_re <= _T_5239_re;
    _T_5240_im <= _T_5239_im;
    _T_5241_re <= _T_5240_re;
    _T_5241_im <= _T_5240_im;
    _T_5242_re <= _T_5241_re;
    _T_5242_im <= _T_5241_im;
    _T_5243_re <= _T_5242_re;
    _T_5243_im <= _T_5242_im;
    _T_5244_re <= _T_5243_re;
    _T_5244_im <= _T_5243_im;
    _T_5245_re <= _T_5244_re;
    _T_5245_im <= _T_5244_im;
    _T_5246_re <= _T_5245_re;
    _T_5246_im <= _T_5245_im;
    _T_5247_re <= _T_5246_re;
    _T_5247_im <= _T_5246_im;
    _T_5248_re <= _T_5247_re;
    _T_5248_im <= _T_5247_im;
    _T_5249_re <= _T_5248_re;
    _T_5249_im <= _T_5248_im;
    _T_5250_re <= _T_5249_re;
    _T_5250_im <= _T_5249_im;
    _T_5251_re <= _T_5250_re;
    _T_5251_im <= _T_5250_im;
    _T_5252_re <= _T_5251_re;
    _T_5252_im <= _T_5251_im;
    _T_5253_re <= _T_5252_re;
    _T_5253_im <= _T_5252_im;
    _T_5254_re <= _T_5253_re;
    _T_5254_im <= _T_5253_im;
    _T_5255_re <= _T_5254_re;
    _T_5255_im <= _T_5254_im;
    _T_5256_re <= _T_5255_re;
    _T_5256_im <= _T_5255_im;
    _T_5257_re <= _T_5256_re;
    _T_5257_im <= _T_5256_im;
    _T_5258_re <= _T_5257_re;
    _T_5258_im <= _T_5257_im;
    _T_5259_re <= _T_5258_re;
    _T_5259_im <= _T_5258_im;
    _T_5260_re <= _T_5259_re;
    _T_5260_im <= _T_5259_im;
    _T_5261_re <= _T_5260_re;
    _T_5261_im <= _T_5260_im;
    _T_5262_re <= _T_5261_re;
    _T_5262_im <= _T_5261_im;
    _T_5263_re <= _T_5262_re;
    _T_5263_im <= _T_5262_im;
    _T_5264_re <= _T_5263_re;
    _T_5264_im <= _T_5263_im;
    _T_5265_re <= _T_5264_re;
    _T_5265_im <= _T_5264_im;
    _T_5266_re <= _T_5265_re;
    _T_5266_im <= _T_5265_im;
    _T_5267_re <= _T_5266_re;
    _T_5267_im <= _T_5266_im;
    _T_5268_re <= _T_5267_re;
    _T_5268_im <= _T_5267_im;
    _T_5269_re <= _T_5268_re;
    _T_5269_im <= _T_5268_im;
    _T_5270_re <= _T_5269_re;
    _T_5270_im <= _T_5269_im;
    _T_5271_re <= _T_5270_re;
    _T_5271_im <= _T_5270_im;
    _T_5272_re <= _T_5271_re;
    _T_5272_im <= _T_5271_im;
    _T_5273_re <= _T_5272_re;
    _T_5273_im <= _T_5272_im;
    _T_5274_re <= _T_5273_re;
    _T_5274_im <= _T_5273_im;
    _T_5275_re <= _T_5274_re;
    _T_5275_im <= _T_5274_im;
    _T_5276_re <= _T_5275_re;
    _T_5276_im <= _T_5275_im;
    _T_5277_re <= _T_5276_re;
    _T_5277_im <= _T_5276_im;
    _T_5278_re <= _T_5277_re;
    _T_5278_im <= _T_5277_im;
    _T_5279_re <= _T_5278_re;
    _T_5279_im <= _T_5278_im;
    _T_5280_re <= _T_5279_re;
    _T_5280_im <= _T_5279_im;
    _T_5281_re <= _T_5280_re;
    _T_5281_im <= _T_5280_im;
    _T_5282_re <= _T_5281_re;
    _T_5282_im <= _T_5281_im;
    _T_5283_re <= _T_5282_re;
    _T_5283_im <= _T_5282_im;
    _T_5284_re <= _T_5283_re;
    _T_5284_im <= _T_5283_im;
    _T_5285_re <= _T_5284_re;
    _T_5285_im <= _T_5284_im;
    _T_5286_re <= _T_5285_re;
    _T_5286_im <= _T_5285_im;
    _T_5287_re <= _T_5286_re;
    _T_5287_im <= _T_5286_im;
    _T_5288_re <= _T_5287_re;
    _T_5288_im <= _T_5287_im;
    _T_5289_re <= _T_5288_re;
    _T_5289_im <= _T_5288_im;
    _T_5290_re <= _T_5289_re;
    _T_5290_im <= _T_5289_im;
    _T_5291_re <= _T_5290_re;
    _T_5291_im <= _T_5290_im;
    _T_5292_re <= _T_5291_re;
    _T_5292_im <= _T_5291_im;
    _T_5293_re <= _T_5292_re;
    _T_5293_im <= _T_5292_im;
    _T_5294_re <= _T_5293_re;
    _T_5294_im <= _T_5293_im;
    _T_5295_re <= _T_5294_re;
    _T_5295_im <= _T_5294_im;
    _T_5296_re <= _T_5295_re;
    _T_5296_im <= _T_5295_im;
    _T_5297_re <= _T_5296_re;
    _T_5297_im <= _T_5296_im;
    _T_5298_re <= _T_5297_re;
    _T_5298_im <= _T_5297_im;
    _T_5299_re <= _T_5298_re;
    _T_5299_im <= _T_5298_im;
    _T_5300_re <= _T_5299_re;
    _T_5300_im <= _T_5299_im;
    _T_5301_re <= _T_5300_re;
    _T_5301_im <= _T_5300_im;
    _T_5302_re <= _T_5301_re;
    _T_5302_im <= _T_5301_im;
    _T_5303_re <= _T_5302_re;
    _T_5303_im <= _T_5302_im;
    _T_5304_re <= _T_5303_re;
    _T_5304_im <= _T_5303_im;
    _T_5305_re <= _T_5304_re;
    _T_5305_im <= _T_5304_im;
    _T_5306_re <= _T_5305_re;
    _T_5306_im <= _T_5305_im;
    _T_5307_re <= _T_5306_re;
    _T_5307_im <= _T_5306_im;
    _T_5308_re <= _T_5307_re;
    _T_5308_im <= _T_5307_im;
    _T_5309_re <= _T_5308_re;
    _T_5309_im <= _T_5308_im;
    _T_5310_re <= _T_5309_re;
    _T_5310_im <= _T_5309_im;
    _T_5311_re <= _T_5310_re;
    _T_5311_im <= _T_5310_im;
    _T_5312_re <= _T_5311_re;
    _T_5312_im <= _T_5311_im;
    _T_5313_re <= _T_5312_re;
    _T_5313_im <= _T_5312_im;
    _T_5314_re <= _T_5313_re;
    _T_5314_im <= _T_5313_im;
    _T_5315_re <= _T_5314_re;
    _T_5315_im <= _T_5314_im;
    _T_5316_re <= _T_5315_re;
    _T_5316_im <= _T_5315_im;
    _T_5317_re <= _T_5316_re;
    _T_5317_im <= _T_5316_im;
    _T_5318_re <= _T_5317_re;
    _T_5318_im <= _T_5317_im;
    _T_5319_re <= _T_5318_re;
    _T_5319_im <= _T_5318_im;
    _T_5320_re <= _T_5319_re;
    _T_5320_im <= _T_5319_im;
    _T_5321_re <= _T_5320_re;
    _T_5321_im <= _T_5320_im;
    _T_5322_re <= _T_5321_re;
    _T_5322_im <= _T_5321_im;
    _T_5325_re <= Butterfly_2_io_out2_re;
    _T_5325_im <= Butterfly_2_io_out2_im;
    _T_5326_re <= _T_5325_re;
    _T_5326_im <= _T_5325_im;
    _T_5327_re <= _T_5326_re;
    _T_5327_im <= _T_5326_im;
    _T_5328_re <= _T_5327_re;
    _T_5328_im <= _T_5327_im;
    _T_5329_re <= _T_5328_re;
    _T_5329_im <= _T_5328_im;
    _T_5330_re <= _T_5329_re;
    _T_5330_im <= _T_5329_im;
    _T_5331_re <= _T_5330_re;
    _T_5331_im <= _T_5330_im;
    _T_5332_re <= _T_5331_re;
    _T_5332_im <= _T_5331_im;
    _T_5333_re <= _T_5332_re;
    _T_5333_im <= _T_5332_im;
    _T_5334_re <= _T_5333_re;
    _T_5334_im <= _T_5333_im;
    _T_5335_re <= _T_5334_re;
    _T_5335_im <= _T_5334_im;
    _T_5336_re <= _T_5335_re;
    _T_5336_im <= _T_5335_im;
    _T_5337_re <= _T_5336_re;
    _T_5337_im <= _T_5336_im;
    _T_5338_re <= _T_5337_re;
    _T_5338_im <= _T_5337_im;
    _T_5339_re <= _T_5338_re;
    _T_5339_im <= _T_5338_im;
    _T_5340_re <= _T_5339_re;
    _T_5340_im <= _T_5339_im;
    _T_5341_re <= _T_5340_re;
    _T_5341_im <= _T_5340_im;
    _T_5342_re <= _T_5341_re;
    _T_5342_im <= _T_5341_im;
    _T_5343_re <= _T_5342_re;
    _T_5343_im <= _T_5342_im;
    _T_5344_re <= _T_5343_re;
    _T_5344_im <= _T_5343_im;
    _T_5345_re <= _T_5344_re;
    _T_5345_im <= _T_5344_im;
    _T_5346_re <= _T_5345_re;
    _T_5346_im <= _T_5345_im;
    _T_5347_re <= _T_5346_re;
    _T_5347_im <= _T_5346_im;
    _T_5348_re <= _T_5347_re;
    _T_5348_im <= _T_5347_im;
    _T_5349_re <= _T_5348_re;
    _T_5349_im <= _T_5348_im;
    _T_5350_re <= _T_5349_re;
    _T_5350_im <= _T_5349_im;
    _T_5351_re <= _T_5350_re;
    _T_5351_im <= _T_5350_im;
    _T_5352_re <= _T_5351_re;
    _T_5352_im <= _T_5351_im;
    _T_5353_re <= _T_5352_re;
    _T_5353_im <= _T_5352_im;
    _T_5354_re <= _T_5353_re;
    _T_5354_im <= _T_5353_im;
    _T_5355_re <= _T_5354_re;
    _T_5355_im <= _T_5354_im;
    _T_5356_re <= _T_5355_re;
    _T_5356_im <= _T_5355_im;
    _T_5357_re <= _T_5356_re;
    _T_5357_im <= _T_5356_im;
    _T_5358_re <= _T_5357_re;
    _T_5358_im <= _T_5357_im;
    _T_5359_re <= _T_5358_re;
    _T_5359_im <= _T_5358_im;
    _T_5360_re <= _T_5359_re;
    _T_5360_im <= _T_5359_im;
    _T_5361_re <= _T_5360_re;
    _T_5361_im <= _T_5360_im;
    _T_5362_re <= _T_5361_re;
    _T_5362_im <= _T_5361_im;
    _T_5363_re <= _T_5362_re;
    _T_5363_im <= _T_5362_im;
    _T_5364_re <= _T_5363_re;
    _T_5364_im <= _T_5363_im;
    _T_5365_re <= _T_5364_re;
    _T_5365_im <= _T_5364_im;
    _T_5366_re <= _T_5365_re;
    _T_5366_im <= _T_5365_im;
    _T_5367_re <= _T_5366_re;
    _T_5367_im <= _T_5366_im;
    _T_5368_re <= _T_5367_re;
    _T_5368_im <= _T_5367_im;
    _T_5369_re <= _T_5368_re;
    _T_5369_im <= _T_5368_im;
    _T_5370_re <= _T_5369_re;
    _T_5370_im <= _T_5369_im;
    _T_5371_re <= _T_5370_re;
    _T_5371_im <= _T_5370_im;
    _T_5372_re <= _T_5371_re;
    _T_5372_im <= _T_5371_im;
    _T_5373_re <= _T_5372_re;
    _T_5373_im <= _T_5372_im;
    _T_5374_re <= _T_5373_re;
    _T_5374_im <= _T_5373_im;
    _T_5375_re <= _T_5374_re;
    _T_5375_im <= _T_5374_im;
    _T_5376_re <= _T_5375_re;
    _T_5376_im <= _T_5375_im;
    _T_5377_re <= _T_5376_re;
    _T_5377_im <= _T_5376_im;
    _T_5378_re <= _T_5377_re;
    _T_5378_im <= _T_5377_im;
    _T_5379_re <= _T_5378_re;
    _T_5379_im <= _T_5378_im;
    _T_5380_re <= _T_5379_re;
    _T_5380_im <= _T_5379_im;
    _T_5381_re <= _T_5380_re;
    _T_5381_im <= _T_5380_im;
    _T_5382_re <= _T_5381_re;
    _T_5382_im <= _T_5381_im;
    _T_5383_re <= _T_5382_re;
    _T_5383_im <= _T_5382_im;
    _T_5384_re <= _T_5383_re;
    _T_5384_im <= _T_5383_im;
    _T_5385_re <= _T_5384_re;
    _T_5385_im <= _T_5384_im;
    _T_5386_re <= _T_5385_re;
    _T_5386_im <= _T_5385_im;
    _T_5387_re <= _T_5386_re;
    _T_5387_im <= _T_5386_im;
    _T_5388_re <= _T_5387_re;
    _T_5388_im <= _T_5387_im;
    _T_5389_re <= _T_5388_re;
    _T_5389_im <= _T_5388_im;
    _T_5390_re <= _T_5389_re;
    _T_5390_im <= _T_5389_im;
    _T_5391_re <= _T_5390_re;
    _T_5391_im <= _T_5390_im;
    _T_5392_re <= _T_5391_re;
    _T_5392_im <= _T_5391_im;
    _T_5393_re <= _T_5392_re;
    _T_5393_im <= _T_5392_im;
    _T_5394_re <= _T_5393_re;
    _T_5394_im <= _T_5393_im;
    _T_5395_re <= _T_5394_re;
    _T_5395_im <= _T_5394_im;
    _T_5396_re <= _T_5395_re;
    _T_5396_im <= _T_5395_im;
    _T_5397_re <= _T_5396_re;
    _T_5397_im <= _T_5396_im;
    _T_5398_re <= _T_5397_re;
    _T_5398_im <= _T_5397_im;
    _T_5399_re <= _T_5398_re;
    _T_5399_im <= _T_5398_im;
    _T_5400_re <= _T_5399_re;
    _T_5400_im <= _T_5399_im;
    _T_5401_re <= _T_5400_re;
    _T_5401_im <= _T_5400_im;
    _T_5402_re <= _T_5401_re;
    _T_5402_im <= _T_5401_im;
    _T_5403_re <= _T_5402_re;
    _T_5403_im <= _T_5402_im;
    _T_5404_re <= _T_5403_re;
    _T_5404_im <= _T_5403_im;
    _T_5405_re <= _T_5404_re;
    _T_5405_im <= _T_5404_im;
    _T_5406_re <= _T_5405_re;
    _T_5406_im <= _T_5405_im;
    _T_5407_re <= _T_5406_re;
    _T_5407_im <= _T_5406_im;
    _T_5408_re <= _T_5407_re;
    _T_5408_im <= _T_5407_im;
    _T_5409_re <= _T_5408_re;
    _T_5409_im <= _T_5408_im;
    _T_5410_re <= _T_5409_re;
    _T_5410_im <= _T_5409_im;
    _T_5411_re <= _T_5410_re;
    _T_5411_im <= _T_5410_im;
    _T_5412_re <= _T_5411_re;
    _T_5412_im <= _T_5411_im;
    _T_5413_re <= _T_5412_re;
    _T_5413_im <= _T_5412_im;
    _T_5414_re <= _T_5413_re;
    _T_5414_im <= _T_5413_im;
    _T_5415_re <= _T_5414_re;
    _T_5415_im <= _T_5414_im;
    _T_5416_re <= _T_5415_re;
    _T_5416_im <= _T_5415_im;
    _T_5417_re <= _T_5416_re;
    _T_5417_im <= _T_5416_im;
    _T_5418_re <= _T_5417_re;
    _T_5418_im <= _T_5417_im;
    _T_5419_re <= _T_5418_re;
    _T_5419_im <= _T_5418_im;
    _T_5420_re <= _T_5419_re;
    _T_5420_im <= _T_5419_im;
    _T_5421_re <= _T_5420_re;
    _T_5421_im <= _T_5420_im;
    _T_5422_re <= _T_5421_re;
    _T_5422_im <= _T_5421_im;
    _T_5423_re <= _T_5422_re;
    _T_5423_im <= _T_5422_im;
    _T_5424_re <= _T_5423_re;
    _T_5424_im <= _T_5423_im;
    _T_5425_re <= _T_5424_re;
    _T_5425_im <= _T_5424_im;
    _T_5426_re <= _T_5425_re;
    _T_5426_im <= _T_5425_im;
    _T_5427_re <= _T_5426_re;
    _T_5427_im <= _T_5426_im;
    _T_5428_re <= _T_5427_re;
    _T_5428_im <= _T_5427_im;
    _T_5429_re <= _T_5428_re;
    _T_5429_im <= _T_5428_im;
    _T_5430_re <= _T_5429_re;
    _T_5430_im <= _T_5429_im;
    _T_5431_re <= _T_5430_re;
    _T_5431_im <= _T_5430_im;
    _T_5432_re <= _T_5431_re;
    _T_5432_im <= _T_5431_im;
    _T_5433_re <= _T_5432_re;
    _T_5433_im <= _T_5432_im;
    _T_5434_re <= _T_5433_re;
    _T_5434_im <= _T_5433_im;
    _T_5435_re <= _T_5434_re;
    _T_5435_im <= _T_5434_im;
    _T_5436_re <= _T_5435_re;
    _T_5436_im <= _T_5435_im;
    _T_5437_re <= _T_5436_re;
    _T_5437_im <= _T_5436_im;
    _T_5438_re <= _T_5437_re;
    _T_5438_im <= _T_5437_im;
    _T_5439_re <= _T_5438_re;
    _T_5439_im <= _T_5438_im;
    _T_5440_re <= _T_5439_re;
    _T_5440_im <= _T_5439_im;
    _T_5441_re <= _T_5440_re;
    _T_5441_im <= _T_5440_im;
    _T_5442_re <= _T_5441_re;
    _T_5442_im <= _T_5441_im;
    _T_5443_re <= _T_5442_re;
    _T_5443_im <= _T_5442_im;
    _T_5444_re <= _T_5443_re;
    _T_5444_im <= _T_5443_im;
    _T_5445_re <= _T_5444_re;
    _T_5445_im <= _T_5444_im;
    _T_5446_re <= _T_5445_re;
    _T_5446_im <= _T_5445_im;
    _T_5447_re <= _T_5446_re;
    _T_5447_im <= _T_5446_im;
    _T_5448_re <= _T_5447_re;
    _T_5448_im <= _T_5447_im;
    _T_5449_re <= _T_5448_re;
    _T_5449_im <= _T_5448_im;
    _T_5450_re <= _T_5449_re;
    _T_5450_im <= _T_5449_im;
    _T_5451_re <= _T_5450_re;
    _T_5451_im <= _T_5450_im;
    _T_5452_re <= _T_5451_re;
    _T_5452_im <= _T_5451_im;
    _T_5453_re <= _T_5452_re;
    _T_5453_im <= _T_5452_im;
    _T_5454_re <= _T_5453_re;
    _T_5454_im <= _T_5453_im;
    _T_5455_re <= _T_5454_re;
    _T_5455_im <= _T_5454_im;
    _T_5456_re <= _T_5455_re;
    _T_5456_im <= _T_5455_im;
    _T_5457_re <= _T_5456_re;
    _T_5457_im <= _T_5456_im;
    _T_5458_re <= _T_5457_re;
    _T_5458_im <= _T_5457_im;
    _T_5459_re <= _T_5458_re;
    _T_5459_im <= _T_5458_im;
    _T_5460_re <= _T_5459_re;
    _T_5460_im <= _T_5459_im;
    _T_5461_re <= _T_5460_re;
    _T_5461_im <= _T_5460_im;
    _T_5462_re <= _T_5461_re;
    _T_5462_im <= _T_5461_im;
    _T_5463_re <= _T_5462_re;
    _T_5463_im <= _T_5462_im;
    _T_5464_re <= _T_5463_re;
    _T_5464_im <= _T_5463_im;
    _T_5465_re <= _T_5464_re;
    _T_5465_im <= _T_5464_im;
    _T_5466_re <= _T_5465_re;
    _T_5466_im <= _T_5465_im;
    _T_5467_re <= _T_5466_re;
    _T_5467_im <= _T_5466_im;
    _T_5468_re <= _T_5467_re;
    _T_5468_im <= _T_5467_im;
    _T_5469_re <= _T_5468_re;
    _T_5469_im <= _T_5468_im;
    _T_5470_re <= _T_5469_re;
    _T_5470_im <= _T_5469_im;
    _T_5471_re <= _T_5470_re;
    _T_5471_im <= _T_5470_im;
    _T_5472_re <= _T_5471_re;
    _T_5472_im <= _T_5471_im;
    _T_5473_re <= _T_5472_re;
    _T_5473_im <= _T_5472_im;
    _T_5474_re <= _T_5473_re;
    _T_5474_im <= _T_5473_im;
    _T_5475_re <= _T_5474_re;
    _T_5475_im <= _T_5474_im;
    _T_5476_re <= _T_5475_re;
    _T_5476_im <= _T_5475_im;
    _T_5477_re <= _T_5476_re;
    _T_5477_im <= _T_5476_im;
    _T_5478_re <= _T_5477_re;
    _T_5478_im <= _T_5477_im;
    _T_5479_re <= _T_5478_re;
    _T_5479_im <= _T_5478_im;
    _T_5480_re <= _T_5479_re;
    _T_5480_im <= _T_5479_im;
    _T_5481_re <= _T_5480_re;
    _T_5481_im <= _T_5480_im;
    _T_5482_re <= _T_5481_re;
    _T_5482_im <= _T_5481_im;
    _T_5483_re <= _T_5482_re;
    _T_5483_im <= _T_5482_im;
    _T_5484_re <= _T_5483_re;
    _T_5484_im <= _T_5483_im;
    _T_5485_re <= _T_5484_re;
    _T_5485_im <= _T_5484_im;
    _T_5486_re <= _T_5485_re;
    _T_5486_im <= _T_5485_im;
    _T_5487_re <= _T_5486_re;
    _T_5487_im <= _T_5486_im;
    _T_5488_re <= _T_5487_re;
    _T_5488_im <= _T_5487_im;
    _T_5489_re <= _T_5488_re;
    _T_5489_im <= _T_5488_im;
    _T_5490_re <= _T_5489_re;
    _T_5490_im <= _T_5489_im;
    _T_5491_re <= _T_5490_re;
    _T_5491_im <= _T_5490_im;
    _T_5492_re <= _T_5491_re;
    _T_5492_im <= _T_5491_im;
    _T_5493_re <= _T_5492_re;
    _T_5493_im <= _T_5492_im;
    _T_5494_re <= _T_5493_re;
    _T_5494_im <= _T_5493_im;
    _T_5495_re <= _T_5494_re;
    _T_5495_im <= _T_5494_im;
    _T_5496_re <= _T_5495_re;
    _T_5496_im <= _T_5495_im;
    _T_5497_re <= _T_5496_re;
    _T_5497_im <= _T_5496_im;
    _T_5498_re <= _T_5497_re;
    _T_5498_im <= _T_5497_im;
    _T_5499_re <= _T_5498_re;
    _T_5499_im <= _T_5498_im;
    _T_5500_re <= _T_5499_re;
    _T_5500_im <= _T_5499_im;
    _T_5501_re <= _T_5500_re;
    _T_5501_im <= _T_5500_im;
    _T_5502_re <= _T_5501_re;
    _T_5502_im <= _T_5501_im;
    _T_5503_re <= _T_5502_re;
    _T_5503_im <= _T_5502_im;
    _T_5504_re <= _T_5503_re;
    _T_5504_im <= _T_5503_im;
    _T_5505_re <= _T_5504_re;
    _T_5505_im <= _T_5504_im;
    _T_5506_re <= _T_5505_re;
    _T_5506_im <= _T_5505_im;
    _T_5507_re <= _T_5506_re;
    _T_5507_im <= _T_5506_im;
    _T_5508_re <= _T_5507_re;
    _T_5508_im <= _T_5507_im;
    _T_5509_re <= _T_5508_re;
    _T_5509_im <= _T_5508_im;
    _T_5510_re <= _T_5509_re;
    _T_5510_im <= _T_5509_im;
    _T_5511_re <= _T_5510_re;
    _T_5511_im <= _T_5510_im;
    _T_5512_re <= _T_5511_re;
    _T_5512_im <= _T_5511_im;
    _T_5513_re <= _T_5512_re;
    _T_5513_im <= _T_5512_im;
    _T_5514_re <= _T_5513_re;
    _T_5514_im <= _T_5513_im;
    _T_5515_re <= _T_5514_re;
    _T_5515_im <= _T_5514_im;
    _T_5516_re <= _T_5515_re;
    _T_5516_im <= _T_5515_im;
    _T_5517_re <= _T_5516_re;
    _T_5517_im <= _T_5516_im;
    _T_5518_re <= _T_5517_re;
    _T_5518_im <= _T_5517_im;
    _T_5519_re <= _T_5518_re;
    _T_5519_im <= _T_5518_im;
    _T_5520_re <= _T_5519_re;
    _T_5520_im <= _T_5519_im;
    _T_5521_re <= _T_5520_re;
    _T_5521_im <= _T_5520_im;
    _T_5522_re <= _T_5521_re;
    _T_5522_im <= _T_5521_im;
    _T_5523_re <= _T_5522_re;
    _T_5523_im <= _T_5522_im;
    _T_5524_re <= _T_5523_re;
    _T_5524_im <= _T_5523_im;
    _T_5525_re <= _T_5524_re;
    _T_5525_im <= _T_5524_im;
    _T_5526_re <= _T_5525_re;
    _T_5526_im <= _T_5525_im;
    _T_5527_re <= _T_5526_re;
    _T_5527_im <= _T_5526_im;
    _T_5528_re <= _T_5527_re;
    _T_5528_im <= _T_5527_im;
    _T_5529_re <= _T_5528_re;
    _T_5529_im <= _T_5528_im;
    _T_5530_re <= _T_5529_re;
    _T_5530_im <= _T_5529_im;
    _T_5531_re <= _T_5530_re;
    _T_5531_im <= _T_5530_im;
    _T_5532_re <= _T_5531_re;
    _T_5532_im <= _T_5531_im;
    _T_5533_re <= _T_5532_re;
    _T_5533_im <= _T_5532_im;
    _T_5534_re <= _T_5533_re;
    _T_5534_im <= _T_5533_im;
    _T_5535_re <= _T_5534_re;
    _T_5535_im <= _T_5534_im;
    _T_5536_re <= _T_5535_re;
    _T_5536_im <= _T_5535_im;
    _T_5537_re <= _T_5536_re;
    _T_5537_im <= _T_5536_im;
    _T_5538_re <= _T_5537_re;
    _T_5538_im <= _T_5537_im;
    _T_5539_re <= _T_5538_re;
    _T_5539_im <= _T_5538_im;
    _T_5540_re <= _T_5539_re;
    _T_5540_im <= _T_5539_im;
    _T_5541_re <= _T_5540_re;
    _T_5541_im <= _T_5540_im;
    _T_5542_re <= _T_5541_re;
    _T_5542_im <= _T_5541_im;
    _T_5543_re <= _T_5542_re;
    _T_5543_im <= _T_5542_im;
    _T_5544_re <= _T_5543_re;
    _T_5544_im <= _T_5543_im;
    _T_5545_re <= _T_5544_re;
    _T_5545_im <= _T_5544_im;
    _T_5546_re <= _T_5545_re;
    _T_5546_im <= _T_5545_im;
    _T_5547_re <= _T_5546_re;
    _T_5547_im <= _T_5546_im;
    _T_5548_re <= _T_5547_re;
    _T_5548_im <= _T_5547_im;
    _T_5549_re <= _T_5548_re;
    _T_5549_im <= _T_5548_im;
    _T_5550_re <= _T_5549_re;
    _T_5550_im <= _T_5549_im;
    _T_5551_re <= _T_5550_re;
    _T_5551_im <= _T_5550_im;
    _T_5552_re <= _T_5551_re;
    _T_5552_im <= _T_5551_im;
    _T_5553_re <= _T_5552_re;
    _T_5553_im <= _T_5552_im;
    _T_5554_re <= _T_5553_re;
    _T_5554_im <= _T_5553_im;
    _T_5555_re <= _T_5554_re;
    _T_5555_im <= _T_5554_im;
    _T_5556_re <= _T_5555_re;
    _T_5556_im <= _T_5555_im;
    _T_5557_re <= _T_5556_re;
    _T_5557_im <= _T_5556_im;
    _T_5558_re <= _T_5557_re;
    _T_5558_im <= _T_5557_im;
    _T_5559_re <= _T_5558_re;
    _T_5559_im <= _T_5558_im;
    _T_5560_re <= _T_5559_re;
    _T_5560_im <= _T_5559_im;
    _T_5561_re <= _T_5560_re;
    _T_5561_im <= _T_5560_im;
    _T_5562_re <= _T_5561_re;
    _T_5562_im <= _T_5561_im;
    _T_5563_re <= _T_5562_re;
    _T_5563_im <= _T_5562_im;
    _T_5564_re <= _T_5563_re;
    _T_5564_im <= _T_5563_im;
    _T_5565_re <= _T_5564_re;
    _T_5565_im <= _T_5564_im;
    _T_5566_re <= _T_5565_re;
    _T_5566_im <= _T_5565_im;
    _T_5567_re <= _T_5566_re;
    _T_5567_im <= _T_5566_im;
    _T_5568_re <= _T_5567_re;
    _T_5568_im <= _T_5567_im;
    _T_5569_re <= _T_5568_re;
    _T_5569_im <= _T_5568_im;
    _T_5570_re <= _T_5569_re;
    _T_5570_im <= _T_5569_im;
    _T_5571_re <= _T_5570_re;
    _T_5571_im <= _T_5570_im;
    _T_5572_re <= _T_5571_re;
    _T_5572_im <= _T_5571_im;
    _T_5573_re <= _T_5572_re;
    _T_5573_im <= _T_5572_im;
    _T_5574_re <= _T_5573_re;
    _T_5574_im <= _T_5573_im;
    _T_5575_re <= _T_5574_re;
    _T_5575_im <= _T_5574_im;
    _T_5576_re <= _T_5575_re;
    _T_5576_im <= _T_5575_im;
    _T_5577_re <= _T_5576_re;
    _T_5577_im <= _T_5576_im;
    _T_5578_re <= _T_5577_re;
    _T_5578_im <= _T_5577_im;
    _T_5579_re <= _T_5578_re;
    _T_5579_im <= _T_5578_im;
    _T_5580_re <= _T_5579_re;
    _T_5580_im <= _T_5579_im;
    _T_5586_re <= Switch_2_io_out1_re;
    _T_5586_im <= Switch_2_io_out1_im;
    _T_5587_re <= _T_5586_re;
    _T_5587_im <= _T_5586_im;
    _T_5588_re <= _T_5587_re;
    _T_5588_im <= _T_5587_im;
    _T_5589_re <= _T_5588_re;
    _T_5589_im <= _T_5588_im;
    _T_5590_re <= _T_5589_re;
    _T_5590_im <= _T_5589_im;
    _T_5591_re <= _T_5590_re;
    _T_5591_im <= _T_5590_im;
    _T_5592_re <= _T_5591_re;
    _T_5592_im <= _T_5591_im;
    _T_5593_re <= _T_5592_re;
    _T_5593_im <= _T_5592_im;
    _T_5594_re <= _T_5593_re;
    _T_5594_im <= _T_5593_im;
    _T_5595_re <= _T_5594_re;
    _T_5595_im <= _T_5594_im;
    _T_5596_re <= _T_5595_re;
    _T_5596_im <= _T_5595_im;
    _T_5597_re <= _T_5596_re;
    _T_5597_im <= _T_5596_im;
    _T_5598_re <= _T_5597_re;
    _T_5598_im <= _T_5597_im;
    _T_5599_re <= _T_5598_re;
    _T_5599_im <= _T_5598_im;
    _T_5600_re <= _T_5599_re;
    _T_5600_im <= _T_5599_im;
    _T_5601_re <= _T_5600_re;
    _T_5601_im <= _T_5600_im;
    _T_5602_re <= _T_5601_re;
    _T_5602_im <= _T_5601_im;
    _T_5603_re <= _T_5602_re;
    _T_5603_im <= _T_5602_im;
    _T_5604_re <= _T_5603_re;
    _T_5604_im <= _T_5603_im;
    _T_5605_re <= _T_5604_re;
    _T_5605_im <= _T_5604_im;
    _T_5606_re <= _T_5605_re;
    _T_5606_im <= _T_5605_im;
    _T_5607_re <= _T_5606_re;
    _T_5607_im <= _T_5606_im;
    _T_5608_re <= _T_5607_re;
    _T_5608_im <= _T_5607_im;
    _T_5609_re <= _T_5608_re;
    _T_5609_im <= _T_5608_im;
    _T_5610_re <= _T_5609_re;
    _T_5610_im <= _T_5609_im;
    _T_5611_re <= _T_5610_re;
    _T_5611_im <= _T_5610_im;
    _T_5612_re <= _T_5611_re;
    _T_5612_im <= _T_5611_im;
    _T_5613_re <= _T_5612_re;
    _T_5613_im <= _T_5612_im;
    _T_5614_re <= _T_5613_re;
    _T_5614_im <= _T_5613_im;
    _T_5615_re <= _T_5614_re;
    _T_5615_im <= _T_5614_im;
    _T_5616_re <= _T_5615_re;
    _T_5616_im <= _T_5615_im;
    _T_5617_re <= _T_5616_re;
    _T_5617_im <= _T_5616_im;
    _T_5618_re <= _T_5617_re;
    _T_5618_im <= _T_5617_im;
    _T_5619_re <= _T_5618_re;
    _T_5619_im <= _T_5618_im;
    _T_5620_re <= _T_5619_re;
    _T_5620_im <= _T_5619_im;
    _T_5621_re <= _T_5620_re;
    _T_5621_im <= _T_5620_im;
    _T_5622_re <= _T_5621_re;
    _T_5622_im <= _T_5621_im;
    _T_5623_re <= _T_5622_re;
    _T_5623_im <= _T_5622_im;
    _T_5624_re <= _T_5623_re;
    _T_5624_im <= _T_5623_im;
    _T_5625_re <= _T_5624_re;
    _T_5625_im <= _T_5624_im;
    _T_5626_re <= _T_5625_re;
    _T_5626_im <= _T_5625_im;
    _T_5627_re <= _T_5626_re;
    _T_5627_im <= _T_5626_im;
    _T_5628_re <= _T_5627_re;
    _T_5628_im <= _T_5627_im;
    _T_5629_re <= _T_5628_re;
    _T_5629_im <= _T_5628_im;
    _T_5630_re <= _T_5629_re;
    _T_5630_im <= _T_5629_im;
    _T_5631_re <= _T_5630_re;
    _T_5631_im <= _T_5630_im;
    _T_5632_re <= _T_5631_re;
    _T_5632_im <= _T_5631_im;
    _T_5633_re <= _T_5632_re;
    _T_5633_im <= _T_5632_im;
    _T_5634_re <= _T_5633_re;
    _T_5634_im <= _T_5633_im;
    _T_5635_re <= _T_5634_re;
    _T_5635_im <= _T_5634_im;
    _T_5636_re <= _T_5635_re;
    _T_5636_im <= _T_5635_im;
    _T_5637_re <= _T_5636_re;
    _T_5637_im <= _T_5636_im;
    _T_5638_re <= _T_5637_re;
    _T_5638_im <= _T_5637_im;
    _T_5639_re <= _T_5638_re;
    _T_5639_im <= _T_5638_im;
    _T_5640_re <= _T_5639_re;
    _T_5640_im <= _T_5639_im;
    _T_5641_re <= _T_5640_re;
    _T_5641_im <= _T_5640_im;
    _T_5642_re <= _T_5641_re;
    _T_5642_im <= _T_5641_im;
    _T_5643_re <= _T_5642_re;
    _T_5643_im <= _T_5642_im;
    _T_5644_re <= _T_5643_re;
    _T_5644_im <= _T_5643_im;
    _T_5645_re <= _T_5644_re;
    _T_5645_im <= _T_5644_im;
    _T_5646_re <= _T_5645_re;
    _T_5646_im <= _T_5645_im;
    _T_5647_re <= _T_5646_re;
    _T_5647_im <= _T_5646_im;
    _T_5648_re <= _T_5647_re;
    _T_5648_im <= _T_5647_im;
    _T_5649_re <= _T_5648_re;
    _T_5649_im <= _T_5648_im;
    _T_5650_re <= _T_5649_re;
    _T_5650_im <= _T_5649_im;
    _T_5651_re <= _T_5650_re;
    _T_5651_im <= _T_5650_im;
    _T_5652_re <= _T_5651_re;
    _T_5652_im <= _T_5651_im;
    _T_5653_re <= _T_5652_re;
    _T_5653_im <= _T_5652_im;
    _T_5654_re <= _T_5653_re;
    _T_5654_im <= _T_5653_im;
    _T_5655_re <= _T_5654_re;
    _T_5655_im <= _T_5654_im;
    _T_5656_re <= _T_5655_re;
    _T_5656_im <= _T_5655_im;
    _T_5657_re <= _T_5656_re;
    _T_5657_im <= _T_5656_im;
    _T_5658_re <= _T_5657_re;
    _T_5658_im <= _T_5657_im;
    _T_5659_re <= _T_5658_re;
    _T_5659_im <= _T_5658_im;
    _T_5660_re <= _T_5659_re;
    _T_5660_im <= _T_5659_im;
    _T_5661_re <= _T_5660_re;
    _T_5661_im <= _T_5660_im;
    _T_5662_re <= _T_5661_re;
    _T_5662_im <= _T_5661_im;
    _T_5663_re <= _T_5662_re;
    _T_5663_im <= _T_5662_im;
    _T_5664_re <= _T_5663_re;
    _T_5664_im <= _T_5663_im;
    _T_5665_re <= _T_5664_re;
    _T_5665_im <= _T_5664_im;
    _T_5666_re <= _T_5665_re;
    _T_5666_im <= _T_5665_im;
    _T_5667_re <= _T_5666_re;
    _T_5667_im <= _T_5666_im;
    _T_5668_re <= _T_5667_re;
    _T_5668_im <= _T_5667_im;
    _T_5669_re <= _T_5668_re;
    _T_5669_im <= _T_5668_im;
    _T_5670_re <= _T_5669_re;
    _T_5670_im <= _T_5669_im;
    _T_5671_re <= _T_5670_re;
    _T_5671_im <= _T_5670_im;
    _T_5672_re <= _T_5671_re;
    _T_5672_im <= _T_5671_im;
    _T_5673_re <= _T_5672_re;
    _T_5673_im <= _T_5672_im;
    _T_5674_re <= _T_5673_re;
    _T_5674_im <= _T_5673_im;
    _T_5675_re <= _T_5674_re;
    _T_5675_im <= _T_5674_im;
    _T_5676_re <= _T_5675_re;
    _T_5676_im <= _T_5675_im;
    _T_5677_re <= _T_5676_re;
    _T_5677_im <= _T_5676_im;
    _T_5678_re <= _T_5677_re;
    _T_5678_im <= _T_5677_im;
    _T_5679_re <= _T_5678_re;
    _T_5679_im <= _T_5678_im;
    _T_5680_re <= _T_5679_re;
    _T_5680_im <= _T_5679_im;
    _T_5681_re <= _T_5680_re;
    _T_5681_im <= _T_5680_im;
    _T_5682_re <= _T_5681_re;
    _T_5682_im <= _T_5681_im;
    _T_5683_re <= _T_5682_re;
    _T_5683_im <= _T_5682_im;
    _T_5684_re <= _T_5683_re;
    _T_5684_im <= _T_5683_im;
    _T_5685_re <= _T_5684_re;
    _T_5685_im <= _T_5684_im;
    _T_5686_re <= _T_5685_re;
    _T_5686_im <= _T_5685_im;
    _T_5687_re <= _T_5686_re;
    _T_5687_im <= _T_5686_im;
    _T_5688_re <= _T_5687_re;
    _T_5688_im <= _T_5687_im;
    _T_5689_re <= _T_5688_re;
    _T_5689_im <= _T_5688_im;
    _T_5690_re <= _T_5689_re;
    _T_5690_im <= _T_5689_im;
    _T_5691_re <= _T_5690_re;
    _T_5691_im <= _T_5690_im;
    _T_5692_re <= _T_5691_re;
    _T_5692_im <= _T_5691_im;
    _T_5693_re <= _T_5692_re;
    _T_5693_im <= _T_5692_im;
    _T_5694_re <= _T_5693_re;
    _T_5694_im <= _T_5693_im;
    _T_5695_re <= _T_5694_re;
    _T_5695_im <= _T_5694_im;
    _T_5696_re <= _T_5695_re;
    _T_5696_im <= _T_5695_im;
    _T_5697_re <= _T_5696_re;
    _T_5697_im <= _T_5696_im;
    _T_5698_re <= _T_5697_re;
    _T_5698_im <= _T_5697_im;
    _T_5699_re <= _T_5698_re;
    _T_5699_im <= _T_5698_im;
    _T_5700_re <= _T_5699_re;
    _T_5700_im <= _T_5699_im;
    _T_5701_re <= _T_5700_re;
    _T_5701_im <= _T_5700_im;
    _T_5702_re <= _T_5701_re;
    _T_5702_im <= _T_5701_im;
    _T_5703_re <= _T_5702_re;
    _T_5703_im <= _T_5702_im;
    _T_5704_re <= _T_5703_re;
    _T_5704_im <= _T_5703_im;
    _T_5705_re <= _T_5704_re;
    _T_5705_im <= _T_5704_im;
    _T_5706_re <= _T_5705_re;
    _T_5706_im <= _T_5705_im;
    _T_5707_re <= _T_5706_re;
    _T_5707_im <= _T_5706_im;
    _T_5708_re <= _T_5707_re;
    _T_5708_im <= _T_5707_im;
    _T_5709_re <= _T_5708_re;
    _T_5709_im <= _T_5708_im;
    _T_5710_re <= _T_5709_re;
    _T_5710_im <= _T_5709_im;
    _T_5711_re <= _T_5710_re;
    _T_5711_im <= _T_5710_im;
    _T_5712_re <= _T_5711_re;
    _T_5712_im <= _T_5711_im;
    _T_5713_re <= _T_5712_re;
    _T_5713_im <= _T_5712_im;
    _T_5714_re <= _T_5713_re;
    _T_5714_im <= _T_5713_im;
    _T_5715_re <= _T_5714_re;
    _T_5715_im <= _T_5714_im;
    _T_5716_re <= _T_5715_re;
    _T_5716_im <= _T_5715_im;
    _T_5717_re <= _T_5716_re;
    _T_5717_im <= _T_5716_im;
    _T_5718_re <= _T_5717_re;
    _T_5718_im <= _T_5717_im;
    _T_5719_re <= _T_5718_re;
    _T_5719_im <= _T_5718_im;
    _T_5720_re <= _T_5719_re;
    _T_5720_im <= _T_5719_im;
    _T_5721_re <= _T_5720_re;
    _T_5721_im <= _T_5720_im;
    _T_5722_re <= _T_5721_re;
    _T_5722_im <= _T_5721_im;
    _T_5723_re <= _T_5722_re;
    _T_5723_im <= _T_5722_im;
    _T_5724_re <= _T_5723_re;
    _T_5724_im <= _T_5723_im;
    _T_5725_re <= _T_5724_re;
    _T_5725_im <= _T_5724_im;
    _T_5726_re <= _T_5725_re;
    _T_5726_im <= _T_5725_im;
    _T_5727_re <= _T_5726_re;
    _T_5727_im <= _T_5726_im;
    _T_5728_re <= _T_5727_re;
    _T_5728_im <= _T_5727_im;
    _T_5729_re <= _T_5728_re;
    _T_5729_im <= _T_5728_im;
    _T_5730_re <= _T_5729_re;
    _T_5730_im <= _T_5729_im;
    _T_5731_re <= _T_5730_re;
    _T_5731_im <= _T_5730_im;
    _T_5732_re <= _T_5731_re;
    _T_5732_im <= _T_5731_im;
    _T_5733_re <= _T_5732_re;
    _T_5733_im <= _T_5732_im;
    _T_5734_re <= _T_5733_re;
    _T_5734_im <= _T_5733_im;
    _T_5735_re <= _T_5734_re;
    _T_5735_im <= _T_5734_im;
    _T_5736_re <= _T_5735_re;
    _T_5736_im <= _T_5735_im;
    _T_5737_re <= _T_5736_re;
    _T_5737_im <= _T_5736_im;
    _T_5738_re <= _T_5737_re;
    _T_5738_im <= _T_5737_im;
    _T_5739_re <= _T_5738_re;
    _T_5739_im <= _T_5738_im;
    _T_5740_re <= _T_5739_re;
    _T_5740_im <= _T_5739_im;
    _T_5741_re <= _T_5740_re;
    _T_5741_im <= _T_5740_im;
    _T_5742_re <= _T_5741_re;
    _T_5742_im <= _T_5741_im;
    _T_5743_re <= _T_5742_re;
    _T_5743_im <= _T_5742_im;
    _T_5744_re <= _T_5743_re;
    _T_5744_im <= _T_5743_im;
    _T_5745_re <= _T_5744_re;
    _T_5745_im <= _T_5744_im;
    _T_5746_re <= _T_5745_re;
    _T_5746_im <= _T_5745_im;
    _T_5747_re <= _T_5746_re;
    _T_5747_im <= _T_5746_im;
    _T_5748_re <= _T_5747_re;
    _T_5748_im <= _T_5747_im;
    _T_5749_re <= _T_5748_re;
    _T_5749_im <= _T_5748_im;
    _T_5750_re <= _T_5749_re;
    _T_5750_im <= _T_5749_im;
    _T_5751_re <= _T_5750_re;
    _T_5751_im <= _T_5750_im;
    _T_5752_re <= _T_5751_re;
    _T_5752_im <= _T_5751_im;
    _T_5753_re <= _T_5752_re;
    _T_5753_im <= _T_5752_im;
    _T_5754_re <= _T_5753_re;
    _T_5754_im <= _T_5753_im;
    _T_5755_re <= _T_5754_re;
    _T_5755_im <= _T_5754_im;
    _T_5756_re <= _T_5755_re;
    _T_5756_im <= _T_5755_im;
    _T_5757_re <= _T_5756_re;
    _T_5757_im <= _T_5756_im;
    _T_5758_re <= _T_5757_re;
    _T_5758_im <= _T_5757_im;
    _T_5759_re <= _T_5758_re;
    _T_5759_im <= _T_5758_im;
    _T_5760_re <= _T_5759_re;
    _T_5760_im <= _T_5759_im;
    _T_5761_re <= _T_5760_re;
    _T_5761_im <= _T_5760_im;
    _T_5762_re <= _T_5761_re;
    _T_5762_im <= _T_5761_im;
    _T_5763_re <= _T_5762_re;
    _T_5763_im <= _T_5762_im;
    _T_5764_re <= _T_5763_re;
    _T_5764_im <= _T_5763_im;
    _T_5765_re <= _T_5764_re;
    _T_5765_im <= _T_5764_im;
    _T_5766_re <= _T_5765_re;
    _T_5766_im <= _T_5765_im;
    _T_5767_re <= _T_5766_re;
    _T_5767_im <= _T_5766_im;
    _T_5768_re <= _T_5767_re;
    _T_5768_im <= _T_5767_im;
    _T_5769_re <= _T_5768_re;
    _T_5769_im <= _T_5768_im;
    _T_5770_re <= _T_5769_re;
    _T_5770_im <= _T_5769_im;
    _T_5771_re <= _T_5770_re;
    _T_5771_im <= _T_5770_im;
    _T_5772_re <= _T_5771_re;
    _T_5772_im <= _T_5771_im;
    _T_5773_re <= _T_5772_re;
    _T_5773_im <= _T_5772_im;
    _T_5774_re <= _T_5773_re;
    _T_5774_im <= _T_5773_im;
    _T_5775_re <= _T_5774_re;
    _T_5775_im <= _T_5774_im;
    _T_5776_re <= _T_5775_re;
    _T_5776_im <= _T_5775_im;
    _T_5777_re <= _T_5776_re;
    _T_5777_im <= _T_5776_im;
    _T_5778_re <= _T_5777_re;
    _T_5778_im <= _T_5777_im;
    _T_5779_re <= _T_5778_re;
    _T_5779_im <= _T_5778_im;
    _T_5780_re <= _T_5779_re;
    _T_5780_im <= _T_5779_im;
    _T_5781_re <= _T_5780_re;
    _T_5781_im <= _T_5780_im;
    _T_5782_re <= _T_5781_re;
    _T_5782_im <= _T_5781_im;
    _T_5783_re <= _T_5782_re;
    _T_5783_im <= _T_5782_im;
    _T_5784_re <= _T_5783_re;
    _T_5784_im <= _T_5783_im;
    _T_5785_re <= _T_5784_re;
    _T_5785_im <= _T_5784_im;
    _T_5786_re <= _T_5785_re;
    _T_5786_im <= _T_5785_im;
    _T_5787_re <= _T_5786_re;
    _T_5787_im <= _T_5786_im;
    _T_5788_re <= _T_5787_re;
    _T_5788_im <= _T_5787_im;
    _T_5789_re <= _T_5788_re;
    _T_5789_im <= _T_5788_im;
    _T_5790_re <= _T_5789_re;
    _T_5790_im <= _T_5789_im;
    _T_5791_re <= _T_5790_re;
    _T_5791_im <= _T_5790_im;
    _T_5792_re <= _T_5791_re;
    _T_5792_im <= _T_5791_im;
    _T_5793_re <= _T_5792_re;
    _T_5793_im <= _T_5792_im;
    _T_5794_re <= _T_5793_re;
    _T_5794_im <= _T_5793_im;
    _T_5795_re <= _T_5794_re;
    _T_5795_im <= _T_5794_im;
    _T_5796_re <= _T_5795_re;
    _T_5796_im <= _T_5795_im;
    _T_5797_re <= _T_5796_re;
    _T_5797_im <= _T_5796_im;
    _T_5798_re <= _T_5797_re;
    _T_5798_im <= _T_5797_im;
    _T_5799_re <= _T_5798_re;
    _T_5799_im <= _T_5798_im;
    _T_5800_re <= _T_5799_re;
    _T_5800_im <= _T_5799_im;
    _T_5801_re <= _T_5800_re;
    _T_5801_im <= _T_5800_im;
    _T_5802_re <= _T_5801_re;
    _T_5802_im <= _T_5801_im;
    _T_5803_re <= _T_5802_re;
    _T_5803_im <= _T_5802_im;
    _T_5804_re <= _T_5803_re;
    _T_5804_im <= _T_5803_im;
    _T_5805_re <= _T_5804_re;
    _T_5805_im <= _T_5804_im;
    _T_5806_re <= _T_5805_re;
    _T_5806_im <= _T_5805_im;
    _T_5807_re <= _T_5806_re;
    _T_5807_im <= _T_5806_im;
    _T_5808_re <= _T_5807_re;
    _T_5808_im <= _T_5807_im;
    _T_5809_re <= _T_5808_re;
    _T_5809_im <= _T_5808_im;
    _T_5810_re <= _T_5809_re;
    _T_5810_im <= _T_5809_im;
    _T_5811_re <= _T_5810_re;
    _T_5811_im <= _T_5810_im;
    _T_5812_re <= _T_5811_re;
    _T_5812_im <= _T_5811_im;
    _T_5813_re <= _T_5812_re;
    _T_5813_im <= _T_5812_im;
    _T_5814_re <= _T_5813_re;
    _T_5814_im <= _T_5813_im;
    _T_5815_re <= _T_5814_re;
    _T_5815_im <= _T_5814_im;
    _T_5816_re <= _T_5815_re;
    _T_5816_im <= _T_5815_im;
    _T_5817_re <= _T_5816_re;
    _T_5817_im <= _T_5816_im;
    _T_5818_re <= _T_5817_re;
    _T_5818_im <= _T_5817_im;
    _T_5819_re <= _T_5818_re;
    _T_5819_im <= _T_5818_im;
    _T_5820_re <= _T_5819_re;
    _T_5820_im <= _T_5819_im;
    _T_5821_re <= _T_5820_re;
    _T_5821_im <= _T_5820_im;
    _T_5822_re <= _T_5821_re;
    _T_5822_im <= _T_5821_im;
    _T_5823_re <= _T_5822_re;
    _T_5823_im <= _T_5822_im;
    _T_5824_re <= _T_5823_re;
    _T_5824_im <= _T_5823_im;
    _T_5825_re <= _T_5824_re;
    _T_5825_im <= _T_5824_im;
    _T_5826_re <= _T_5825_re;
    _T_5826_im <= _T_5825_im;
    _T_5827_re <= _T_5826_re;
    _T_5827_im <= _T_5826_im;
    _T_5828_re <= _T_5827_re;
    _T_5828_im <= _T_5827_im;
    _T_5829_re <= _T_5828_re;
    _T_5829_im <= _T_5828_im;
    _T_5830_re <= _T_5829_re;
    _T_5830_im <= _T_5829_im;
    _T_5831_re <= _T_5830_re;
    _T_5831_im <= _T_5830_im;
    _T_5832_re <= _T_5831_re;
    _T_5832_im <= _T_5831_im;
    _T_5833_re <= _T_5832_re;
    _T_5833_im <= _T_5832_im;
    _T_5834_re <= _T_5833_re;
    _T_5834_im <= _T_5833_im;
    _T_5835_re <= _T_5834_re;
    _T_5835_im <= _T_5834_im;
    _T_5836_re <= _T_5835_re;
    _T_5836_im <= _T_5835_im;
    _T_5837_re <= _T_5836_re;
    _T_5837_im <= _T_5836_im;
    _T_5838_re <= _T_5837_re;
    _T_5838_im <= _T_5837_im;
    _T_5839_re <= _T_5838_re;
    _T_5839_im <= _T_5838_im;
    _T_5840_re <= _T_5839_re;
    _T_5840_im <= _T_5839_im;
    _T_5841_re <= _T_5840_re;
    _T_5841_im <= _T_5840_im;
    _T_5844_re <= Butterfly_3_io_out2_re;
    _T_5844_im <= Butterfly_3_io_out2_im;
    _T_5845_re <= _T_5844_re;
    _T_5845_im <= _T_5844_im;
    _T_5846_re <= _T_5845_re;
    _T_5846_im <= _T_5845_im;
    _T_5847_re <= _T_5846_re;
    _T_5847_im <= _T_5846_im;
    _T_5848_re <= _T_5847_re;
    _T_5848_im <= _T_5847_im;
    _T_5849_re <= _T_5848_re;
    _T_5849_im <= _T_5848_im;
    _T_5850_re <= _T_5849_re;
    _T_5850_im <= _T_5849_im;
    _T_5851_re <= _T_5850_re;
    _T_5851_im <= _T_5850_im;
    _T_5852_re <= _T_5851_re;
    _T_5852_im <= _T_5851_im;
    _T_5853_re <= _T_5852_re;
    _T_5853_im <= _T_5852_im;
    _T_5854_re <= _T_5853_re;
    _T_5854_im <= _T_5853_im;
    _T_5855_re <= _T_5854_re;
    _T_5855_im <= _T_5854_im;
    _T_5856_re <= _T_5855_re;
    _T_5856_im <= _T_5855_im;
    _T_5857_re <= _T_5856_re;
    _T_5857_im <= _T_5856_im;
    _T_5858_re <= _T_5857_re;
    _T_5858_im <= _T_5857_im;
    _T_5859_re <= _T_5858_re;
    _T_5859_im <= _T_5858_im;
    _T_5860_re <= _T_5859_re;
    _T_5860_im <= _T_5859_im;
    _T_5861_re <= _T_5860_re;
    _T_5861_im <= _T_5860_im;
    _T_5862_re <= _T_5861_re;
    _T_5862_im <= _T_5861_im;
    _T_5863_re <= _T_5862_re;
    _T_5863_im <= _T_5862_im;
    _T_5864_re <= _T_5863_re;
    _T_5864_im <= _T_5863_im;
    _T_5865_re <= _T_5864_re;
    _T_5865_im <= _T_5864_im;
    _T_5866_re <= _T_5865_re;
    _T_5866_im <= _T_5865_im;
    _T_5867_re <= _T_5866_re;
    _T_5867_im <= _T_5866_im;
    _T_5868_re <= _T_5867_re;
    _T_5868_im <= _T_5867_im;
    _T_5869_re <= _T_5868_re;
    _T_5869_im <= _T_5868_im;
    _T_5870_re <= _T_5869_re;
    _T_5870_im <= _T_5869_im;
    _T_5871_re <= _T_5870_re;
    _T_5871_im <= _T_5870_im;
    _T_5872_re <= _T_5871_re;
    _T_5872_im <= _T_5871_im;
    _T_5873_re <= _T_5872_re;
    _T_5873_im <= _T_5872_im;
    _T_5874_re <= _T_5873_re;
    _T_5874_im <= _T_5873_im;
    _T_5875_re <= _T_5874_re;
    _T_5875_im <= _T_5874_im;
    _T_5876_re <= _T_5875_re;
    _T_5876_im <= _T_5875_im;
    _T_5877_re <= _T_5876_re;
    _T_5877_im <= _T_5876_im;
    _T_5878_re <= _T_5877_re;
    _T_5878_im <= _T_5877_im;
    _T_5879_re <= _T_5878_re;
    _T_5879_im <= _T_5878_im;
    _T_5880_re <= _T_5879_re;
    _T_5880_im <= _T_5879_im;
    _T_5881_re <= _T_5880_re;
    _T_5881_im <= _T_5880_im;
    _T_5882_re <= _T_5881_re;
    _T_5882_im <= _T_5881_im;
    _T_5883_re <= _T_5882_re;
    _T_5883_im <= _T_5882_im;
    _T_5884_re <= _T_5883_re;
    _T_5884_im <= _T_5883_im;
    _T_5885_re <= _T_5884_re;
    _T_5885_im <= _T_5884_im;
    _T_5886_re <= _T_5885_re;
    _T_5886_im <= _T_5885_im;
    _T_5887_re <= _T_5886_re;
    _T_5887_im <= _T_5886_im;
    _T_5888_re <= _T_5887_re;
    _T_5888_im <= _T_5887_im;
    _T_5889_re <= _T_5888_re;
    _T_5889_im <= _T_5888_im;
    _T_5890_re <= _T_5889_re;
    _T_5890_im <= _T_5889_im;
    _T_5891_re <= _T_5890_re;
    _T_5891_im <= _T_5890_im;
    _T_5892_re <= _T_5891_re;
    _T_5892_im <= _T_5891_im;
    _T_5893_re <= _T_5892_re;
    _T_5893_im <= _T_5892_im;
    _T_5894_re <= _T_5893_re;
    _T_5894_im <= _T_5893_im;
    _T_5895_re <= _T_5894_re;
    _T_5895_im <= _T_5894_im;
    _T_5896_re <= _T_5895_re;
    _T_5896_im <= _T_5895_im;
    _T_5897_re <= _T_5896_re;
    _T_5897_im <= _T_5896_im;
    _T_5898_re <= _T_5897_re;
    _T_5898_im <= _T_5897_im;
    _T_5899_re <= _T_5898_re;
    _T_5899_im <= _T_5898_im;
    _T_5900_re <= _T_5899_re;
    _T_5900_im <= _T_5899_im;
    _T_5901_re <= _T_5900_re;
    _T_5901_im <= _T_5900_im;
    _T_5902_re <= _T_5901_re;
    _T_5902_im <= _T_5901_im;
    _T_5903_re <= _T_5902_re;
    _T_5903_im <= _T_5902_im;
    _T_5904_re <= _T_5903_re;
    _T_5904_im <= _T_5903_im;
    _T_5905_re <= _T_5904_re;
    _T_5905_im <= _T_5904_im;
    _T_5906_re <= _T_5905_re;
    _T_5906_im <= _T_5905_im;
    _T_5907_re <= _T_5906_re;
    _T_5907_im <= _T_5906_im;
    _T_5908_re <= _T_5907_re;
    _T_5908_im <= _T_5907_im;
    _T_5909_re <= _T_5908_re;
    _T_5909_im <= _T_5908_im;
    _T_5910_re <= _T_5909_re;
    _T_5910_im <= _T_5909_im;
    _T_5911_re <= _T_5910_re;
    _T_5911_im <= _T_5910_im;
    _T_5912_re <= _T_5911_re;
    _T_5912_im <= _T_5911_im;
    _T_5913_re <= _T_5912_re;
    _T_5913_im <= _T_5912_im;
    _T_5914_re <= _T_5913_re;
    _T_5914_im <= _T_5913_im;
    _T_5915_re <= _T_5914_re;
    _T_5915_im <= _T_5914_im;
    _T_5916_re <= _T_5915_re;
    _T_5916_im <= _T_5915_im;
    _T_5917_re <= _T_5916_re;
    _T_5917_im <= _T_5916_im;
    _T_5918_re <= _T_5917_re;
    _T_5918_im <= _T_5917_im;
    _T_5919_re <= _T_5918_re;
    _T_5919_im <= _T_5918_im;
    _T_5920_re <= _T_5919_re;
    _T_5920_im <= _T_5919_im;
    _T_5921_re <= _T_5920_re;
    _T_5921_im <= _T_5920_im;
    _T_5922_re <= _T_5921_re;
    _T_5922_im <= _T_5921_im;
    _T_5923_re <= _T_5922_re;
    _T_5923_im <= _T_5922_im;
    _T_5924_re <= _T_5923_re;
    _T_5924_im <= _T_5923_im;
    _T_5925_re <= _T_5924_re;
    _T_5925_im <= _T_5924_im;
    _T_5926_re <= _T_5925_re;
    _T_5926_im <= _T_5925_im;
    _T_5927_re <= _T_5926_re;
    _T_5927_im <= _T_5926_im;
    _T_5928_re <= _T_5927_re;
    _T_5928_im <= _T_5927_im;
    _T_5929_re <= _T_5928_re;
    _T_5929_im <= _T_5928_im;
    _T_5930_re <= _T_5929_re;
    _T_5930_im <= _T_5929_im;
    _T_5931_re <= _T_5930_re;
    _T_5931_im <= _T_5930_im;
    _T_5932_re <= _T_5931_re;
    _T_5932_im <= _T_5931_im;
    _T_5933_re <= _T_5932_re;
    _T_5933_im <= _T_5932_im;
    _T_5934_re <= _T_5933_re;
    _T_5934_im <= _T_5933_im;
    _T_5935_re <= _T_5934_re;
    _T_5935_im <= _T_5934_im;
    _T_5936_re <= _T_5935_re;
    _T_5936_im <= _T_5935_im;
    _T_5937_re <= _T_5936_re;
    _T_5937_im <= _T_5936_im;
    _T_5938_re <= _T_5937_re;
    _T_5938_im <= _T_5937_im;
    _T_5939_re <= _T_5938_re;
    _T_5939_im <= _T_5938_im;
    _T_5940_re <= _T_5939_re;
    _T_5940_im <= _T_5939_im;
    _T_5941_re <= _T_5940_re;
    _T_5941_im <= _T_5940_im;
    _T_5942_re <= _T_5941_re;
    _T_5942_im <= _T_5941_im;
    _T_5943_re <= _T_5942_re;
    _T_5943_im <= _T_5942_im;
    _T_5944_re <= _T_5943_re;
    _T_5944_im <= _T_5943_im;
    _T_5945_re <= _T_5944_re;
    _T_5945_im <= _T_5944_im;
    _T_5946_re <= _T_5945_re;
    _T_5946_im <= _T_5945_im;
    _T_5947_re <= _T_5946_re;
    _T_5947_im <= _T_5946_im;
    _T_5948_re <= _T_5947_re;
    _T_5948_im <= _T_5947_im;
    _T_5949_re <= _T_5948_re;
    _T_5949_im <= _T_5948_im;
    _T_5950_re <= _T_5949_re;
    _T_5950_im <= _T_5949_im;
    _T_5951_re <= _T_5950_re;
    _T_5951_im <= _T_5950_im;
    _T_5952_re <= _T_5951_re;
    _T_5952_im <= _T_5951_im;
    _T_5953_re <= _T_5952_re;
    _T_5953_im <= _T_5952_im;
    _T_5954_re <= _T_5953_re;
    _T_5954_im <= _T_5953_im;
    _T_5955_re <= _T_5954_re;
    _T_5955_im <= _T_5954_im;
    _T_5956_re <= _T_5955_re;
    _T_5956_im <= _T_5955_im;
    _T_5957_re <= _T_5956_re;
    _T_5957_im <= _T_5956_im;
    _T_5958_re <= _T_5957_re;
    _T_5958_im <= _T_5957_im;
    _T_5959_re <= _T_5958_re;
    _T_5959_im <= _T_5958_im;
    _T_5960_re <= _T_5959_re;
    _T_5960_im <= _T_5959_im;
    _T_5961_re <= _T_5960_re;
    _T_5961_im <= _T_5960_im;
    _T_5962_re <= _T_5961_re;
    _T_5962_im <= _T_5961_im;
    _T_5963_re <= _T_5962_re;
    _T_5963_im <= _T_5962_im;
    _T_5964_re <= _T_5963_re;
    _T_5964_im <= _T_5963_im;
    _T_5965_re <= _T_5964_re;
    _T_5965_im <= _T_5964_im;
    _T_5966_re <= _T_5965_re;
    _T_5966_im <= _T_5965_im;
    _T_5967_re <= _T_5966_re;
    _T_5967_im <= _T_5966_im;
    _T_5968_re <= _T_5967_re;
    _T_5968_im <= _T_5967_im;
    _T_5969_re <= _T_5968_re;
    _T_5969_im <= _T_5968_im;
    _T_5970_re <= _T_5969_re;
    _T_5970_im <= _T_5969_im;
    _T_5971_re <= _T_5970_re;
    _T_5971_im <= _T_5970_im;
    _T_5977_re <= Switch_3_io_out1_re;
    _T_5977_im <= Switch_3_io_out1_im;
    _T_5978_re <= _T_5977_re;
    _T_5978_im <= _T_5977_im;
    _T_5979_re <= _T_5978_re;
    _T_5979_im <= _T_5978_im;
    _T_5980_re <= _T_5979_re;
    _T_5980_im <= _T_5979_im;
    _T_5981_re <= _T_5980_re;
    _T_5981_im <= _T_5980_im;
    _T_5982_re <= _T_5981_re;
    _T_5982_im <= _T_5981_im;
    _T_5983_re <= _T_5982_re;
    _T_5983_im <= _T_5982_im;
    _T_5984_re <= _T_5983_re;
    _T_5984_im <= _T_5983_im;
    _T_5985_re <= _T_5984_re;
    _T_5985_im <= _T_5984_im;
    _T_5986_re <= _T_5985_re;
    _T_5986_im <= _T_5985_im;
    _T_5987_re <= _T_5986_re;
    _T_5987_im <= _T_5986_im;
    _T_5988_re <= _T_5987_re;
    _T_5988_im <= _T_5987_im;
    _T_5989_re <= _T_5988_re;
    _T_5989_im <= _T_5988_im;
    _T_5990_re <= _T_5989_re;
    _T_5990_im <= _T_5989_im;
    _T_5991_re <= _T_5990_re;
    _T_5991_im <= _T_5990_im;
    _T_5992_re <= _T_5991_re;
    _T_5992_im <= _T_5991_im;
    _T_5993_re <= _T_5992_re;
    _T_5993_im <= _T_5992_im;
    _T_5994_re <= _T_5993_re;
    _T_5994_im <= _T_5993_im;
    _T_5995_re <= _T_5994_re;
    _T_5995_im <= _T_5994_im;
    _T_5996_re <= _T_5995_re;
    _T_5996_im <= _T_5995_im;
    _T_5997_re <= _T_5996_re;
    _T_5997_im <= _T_5996_im;
    _T_5998_re <= _T_5997_re;
    _T_5998_im <= _T_5997_im;
    _T_5999_re <= _T_5998_re;
    _T_5999_im <= _T_5998_im;
    _T_6000_re <= _T_5999_re;
    _T_6000_im <= _T_5999_im;
    _T_6001_re <= _T_6000_re;
    _T_6001_im <= _T_6000_im;
    _T_6002_re <= _T_6001_re;
    _T_6002_im <= _T_6001_im;
    _T_6003_re <= _T_6002_re;
    _T_6003_im <= _T_6002_im;
    _T_6004_re <= _T_6003_re;
    _T_6004_im <= _T_6003_im;
    _T_6005_re <= _T_6004_re;
    _T_6005_im <= _T_6004_im;
    _T_6006_re <= _T_6005_re;
    _T_6006_im <= _T_6005_im;
    _T_6007_re <= _T_6006_re;
    _T_6007_im <= _T_6006_im;
    _T_6008_re <= _T_6007_re;
    _T_6008_im <= _T_6007_im;
    _T_6009_re <= _T_6008_re;
    _T_6009_im <= _T_6008_im;
    _T_6010_re <= _T_6009_re;
    _T_6010_im <= _T_6009_im;
    _T_6011_re <= _T_6010_re;
    _T_6011_im <= _T_6010_im;
    _T_6012_re <= _T_6011_re;
    _T_6012_im <= _T_6011_im;
    _T_6013_re <= _T_6012_re;
    _T_6013_im <= _T_6012_im;
    _T_6014_re <= _T_6013_re;
    _T_6014_im <= _T_6013_im;
    _T_6015_re <= _T_6014_re;
    _T_6015_im <= _T_6014_im;
    _T_6016_re <= _T_6015_re;
    _T_6016_im <= _T_6015_im;
    _T_6017_re <= _T_6016_re;
    _T_6017_im <= _T_6016_im;
    _T_6018_re <= _T_6017_re;
    _T_6018_im <= _T_6017_im;
    _T_6019_re <= _T_6018_re;
    _T_6019_im <= _T_6018_im;
    _T_6020_re <= _T_6019_re;
    _T_6020_im <= _T_6019_im;
    _T_6021_re <= _T_6020_re;
    _T_6021_im <= _T_6020_im;
    _T_6022_re <= _T_6021_re;
    _T_6022_im <= _T_6021_im;
    _T_6023_re <= _T_6022_re;
    _T_6023_im <= _T_6022_im;
    _T_6024_re <= _T_6023_re;
    _T_6024_im <= _T_6023_im;
    _T_6025_re <= _T_6024_re;
    _T_6025_im <= _T_6024_im;
    _T_6026_re <= _T_6025_re;
    _T_6026_im <= _T_6025_im;
    _T_6027_re <= _T_6026_re;
    _T_6027_im <= _T_6026_im;
    _T_6028_re <= _T_6027_re;
    _T_6028_im <= _T_6027_im;
    _T_6029_re <= _T_6028_re;
    _T_6029_im <= _T_6028_im;
    _T_6030_re <= _T_6029_re;
    _T_6030_im <= _T_6029_im;
    _T_6031_re <= _T_6030_re;
    _T_6031_im <= _T_6030_im;
    _T_6032_re <= _T_6031_re;
    _T_6032_im <= _T_6031_im;
    _T_6033_re <= _T_6032_re;
    _T_6033_im <= _T_6032_im;
    _T_6034_re <= _T_6033_re;
    _T_6034_im <= _T_6033_im;
    _T_6035_re <= _T_6034_re;
    _T_6035_im <= _T_6034_im;
    _T_6036_re <= _T_6035_re;
    _T_6036_im <= _T_6035_im;
    _T_6037_re <= _T_6036_re;
    _T_6037_im <= _T_6036_im;
    _T_6038_re <= _T_6037_re;
    _T_6038_im <= _T_6037_im;
    _T_6039_re <= _T_6038_re;
    _T_6039_im <= _T_6038_im;
    _T_6040_re <= _T_6039_re;
    _T_6040_im <= _T_6039_im;
    _T_6041_re <= _T_6040_re;
    _T_6041_im <= _T_6040_im;
    _T_6042_re <= _T_6041_re;
    _T_6042_im <= _T_6041_im;
    _T_6043_re <= _T_6042_re;
    _T_6043_im <= _T_6042_im;
    _T_6044_re <= _T_6043_re;
    _T_6044_im <= _T_6043_im;
    _T_6045_re <= _T_6044_re;
    _T_6045_im <= _T_6044_im;
    _T_6046_re <= _T_6045_re;
    _T_6046_im <= _T_6045_im;
    _T_6047_re <= _T_6046_re;
    _T_6047_im <= _T_6046_im;
    _T_6048_re <= _T_6047_re;
    _T_6048_im <= _T_6047_im;
    _T_6049_re <= _T_6048_re;
    _T_6049_im <= _T_6048_im;
    _T_6050_re <= _T_6049_re;
    _T_6050_im <= _T_6049_im;
    _T_6051_re <= _T_6050_re;
    _T_6051_im <= _T_6050_im;
    _T_6052_re <= _T_6051_re;
    _T_6052_im <= _T_6051_im;
    _T_6053_re <= _T_6052_re;
    _T_6053_im <= _T_6052_im;
    _T_6054_re <= _T_6053_re;
    _T_6054_im <= _T_6053_im;
    _T_6055_re <= _T_6054_re;
    _T_6055_im <= _T_6054_im;
    _T_6056_re <= _T_6055_re;
    _T_6056_im <= _T_6055_im;
    _T_6057_re <= _T_6056_re;
    _T_6057_im <= _T_6056_im;
    _T_6058_re <= _T_6057_re;
    _T_6058_im <= _T_6057_im;
    _T_6059_re <= _T_6058_re;
    _T_6059_im <= _T_6058_im;
    _T_6060_re <= _T_6059_re;
    _T_6060_im <= _T_6059_im;
    _T_6061_re <= _T_6060_re;
    _T_6061_im <= _T_6060_im;
    _T_6062_re <= _T_6061_re;
    _T_6062_im <= _T_6061_im;
    _T_6063_re <= _T_6062_re;
    _T_6063_im <= _T_6062_im;
    _T_6064_re <= _T_6063_re;
    _T_6064_im <= _T_6063_im;
    _T_6065_re <= _T_6064_re;
    _T_6065_im <= _T_6064_im;
    _T_6066_re <= _T_6065_re;
    _T_6066_im <= _T_6065_im;
    _T_6067_re <= _T_6066_re;
    _T_6067_im <= _T_6066_im;
    _T_6068_re <= _T_6067_re;
    _T_6068_im <= _T_6067_im;
    _T_6069_re <= _T_6068_re;
    _T_6069_im <= _T_6068_im;
    _T_6070_re <= _T_6069_re;
    _T_6070_im <= _T_6069_im;
    _T_6071_re <= _T_6070_re;
    _T_6071_im <= _T_6070_im;
    _T_6072_re <= _T_6071_re;
    _T_6072_im <= _T_6071_im;
    _T_6073_re <= _T_6072_re;
    _T_6073_im <= _T_6072_im;
    _T_6074_re <= _T_6073_re;
    _T_6074_im <= _T_6073_im;
    _T_6075_re <= _T_6074_re;
    _T_6075_im <= _T_6074_im;
    _T_6076_re <= _T_6075_re;
    _T_6076_im <= _T_6075_im;
    _T_6077_re <= _T_6076_re;
    _T_6077_im <= _T_6076_im;
    _T_6078_re <= _T_6077_re;
    _T_6078_im <= _T_6077_im;
    _T_6079_re <= _T_6078_re;
    _T_6079_im <= _T_6078_im;
    _T_6080_re <= _T_6079_re;
    _T_6080_im <= _T_6079_im;
    _T_6081_re <= _T_6080_re;
    _T_6081_im <= _T_6080_im;
    _T_6082_re <= _T_6081_re;
    _T_6082_im <= _T_6081_im;
    _T_6083_re <= _T_6082_re;
    _T_6083_im <= _T_6082_im;
    _T_6084_re <= _T_6083_re;
    _T_6084_im <= _T_6083_im;
    _T_6085_re <= _T_6084_re;
    _T_6085_im <= _T_6084_im;
    _T_6086_re <= _T_6085_re;
    _T_6086_im <= _T_6085_im;
    _T_6087_re <= _T_6086_re;
    _T_6087_im <= _T_6086_im;
    _T_6088_re <= _T_6087_re;
    _T_6088_im <= _T_6087_im;
    _T_6089_re <= _T_6088_re;
    _T_6089_im <= _T_6088_im;
    _T_6090_re <= _T_6089_re;
    _T_6090_im <= _T_6089_im;
    _T_6091_re <= _T_6090_re;
    _T_6091_im <= _T_6090_im;
    _T_6092_re <= _T_6091_re;
    _T_6092_im <= _T_6091_im;
    _T_6093_re <= _T_6092_re;
    _T_6093_im <= _T_6092_im;
    _T_6094_re <= _T_6093_re;
    _T_6094_im <= _T_6093_im;
    _T_6095_re <= _T_6094_re;
    _T_6095_im <= _T_6094_im;
    _T_6096_re <= _T_6095_re;
    _T_6096_im <= _T_6095_im;
    _T_6097_re <= _T_6096_re;
    _T_6097_im <= _T_6096_im;
    _T_6098_re <= _T_6097_re;
    _T_6098_im <= _T_6097_im;
    _T_6099_re <= _T_6098_re;
    _T_6099_im <= _T_6098_im;
    _T_6100_re <= _T_6099_re;
    _T_6100_im <= _T_6099_im;
    _T_6101_re <= _T_6100_re;
    _T_6101_im <= _T_6100_im;
    _T_6102_re <= _T_6101_re;
    _T_6102_im <= _T_6101_im;
    _T_6103_re <= _T_6102_re;
    _T_6103_im <= _T_6102_im;
    _T_6104_re <= _T_6103_re;
    _T_6104_im <= _T_6103_im;
    _T_6107_re <= Butterfly_4_io_out2_re;
    _T_6107_im <= Butterfly_4_io_out2_im;
    _T_6108_re <= _T_6107_re;
    _T_6108_im <= _T_6107_im;
    _T_6109_re <= _T_6108_re;
    _T_6109_im <= _T_6108_im;
    _T_6110_re <= _T_6109_re;
    _T_6110_im <= _T_6109_im;
    _T_6111_re <= _T_6110_re;
    _T_6111_im <= _T_6110_im;
    _T_6112_re <= _T_6111_re;
    _T_6112_im <= _T_6111_im;
    _T_6113_re <= _T_6112_re;
    _T_6113_im <= _T_6112_im;
    _T_6114_re <= _T_6113_re;
    _T_6114_im <= _T_6113_im;
    _T_6115_re <= _T_6114_re;
    _T_6115_im <= _T_6114_im;
    _T_6116_re <= _T_6115_re;
    _T_6116_im <= _T_6115_im;
    _T_6117_re <= _T_6116_re;
    _T_6117_im <= _T_6116_im;
    _T_6118_re <= _T_6117_re;
    _T_6118_im <= _T_6117_im;
    _T_6119_re <= _T_6118_re;
    _T_6119_im <= _T_6118_im;
    _T_6120_re <= _T_6119_re;
    _T_6120_im <= _T_6119_im;
    _T_6121_re <= _T_6120_re;
    _T_6121_im <= _T_6120_im;
    _T_6122_re <= _T_6121_re;
    _T_6122_im <= _T_6121_im;
    _T_6123_re <= _T_6122_re;
    _T_6123_im <= _T_6122_im;
    _T_6124_re <= _T_6123_re;
    _T_6124_im <= _T_6123_im;
    _T_6125_re <= _T_6124_re;
    _T_6125_im <= _T_6124_im;
    _T_6126_re <= _T_6125_re;
    _T_6126_im <= _T_6125_im;
    _T_6127_re <= _T_6126_re;
    _T_6127_im <= _T_6126_im;
    _T_6128_re <= _T_6127_re;
    _T_6128_im <= _T_6127_im;
    _T_6129_re <= _T_6128_re;
    _T_6129_im <= _T_6128_im;
    _T_6130_re <= _T_6129_re;
    _T_6130_im <= _T_6129_im;
    _T_6131_re <= _T_6130_re;
    _T_6131_im <= _T_6130_im;
    _T_6132_re <= _T_6131_re;
    _T_6132_im <= _T_6131_im;
    _T_6133_re <= _T_6132_re;
    _T_6133_im <= _T_6132_im;
    _T_6134_re <= _T_6133_re;
    _T_6134_im <= _T_6133_im;
    _T_6135_re <= _T_6134_re;
    _T_6135_im <= _T_6134_im;
    _T_6136_re <= _T_6135_re;
    _T_6136_im <= _T_6135_im;
    _T_6137_re <= _T_6136_re;
    _T_6137_im <= _T_6136_im;
    _T_6138_re <= _T_6137_re;
    _T_6138_im <= _T_6137_im;
    _T_6139_re <= _T_6138_re;
    _T_6139_im <= _T_6138_im;
    _T_6140_re <= _T_6139_re;
    _T_6140_im <= _T_6139_im;
    _T_6141_re <= _T_6140_re;
    _T_6141_im <= _T_6140_im;
    _T_6142_re <= _T_6141_re;
    _T_6142_im <= _T_6141_im;
    _T_6143_re <= _T_6142_re;
    _T_6143_im <= _T_6142_im;
    _T_6144_re <= _T_6143_re;
    _T_6144_im <= _T_6143_im;
    _T_6145_re <= _T_6144_re;
    _T_6145_im <= _T_6144_im;
    _T_6146_re <= _T_6145_re;
    _T_6146_im <= _T_6145_im;
    _T_6147_re <= _T_6146_re;
    _T_6147_im <= _T_6146_im;
    _T_6148_re <= _T_6147_re;
    _T_6148_im <= _T_6147_im;
    _T_6149_re <= _T_6148_re;
    _T_6149_im <= _T_6148_im;
    _T_6150_re <= _T_6149_re;
    _T_6150_im <= _T_6149_im;
    _T_6151_re <= _T_6150_re;
    _T_6151_im <= _T_6150_im;
    _T_6152_re <= _T_6151_re;
    _T_6152_im <= _T_6151_im;
    _T_6153_re <= _T_6152_re;
    _T_6153_im <= _T_6152_im;
    _T_6154_re <= _T_6153_re;
    _T_6154_im <= _T_6153_im;
    _T_6155_re <= _T_6154_re;
    _T_6155_im <= _T_6154_im;
    _T_6156_re <= _T_6155_re;
    _T_6156_im <= _T_6155_im;
    _T_6157_re <= _T_6156_re;
    _T_6157_im <= _T_6156_im;
    _T_6158_re <= _T_6157_re;
    _T_6158_im <= _T_6157_im;
    _T_6159_re <= _T_6158_re;
    _T_6159_im <= _T_6158_im;
    _T_6160_re <= _T_6159_re;
    _T_6160_im <= _T_6159_im;
    _T_6161_re <= _T_6160_re;
    _T_6161_im <= _T_6160_im;
    _T_6162_re <= _T_6161_re;
    _T_6162_im <= _T_6161_im;
    _T_6163_re <= _T_6162_re;
    _T_6163_im <= _T_6162_im;
    _T_6164_re <= _T_6163_re;
    _T_6164_im <= _T_6163_im;
    _T_6165_re <= _T_6164_re;
    _T_6165_im <= _T_6164_im;
    _T_6166_re <= _T_6165_re;
    _T_6166_im <= _T_6165_im;
    _T_6167_re <= _T_6166_re;
    _T_6167_im <= _T_6166_im;
    _T_6168_re <= _T_6167_re;
    _T_6168_im <= _T_6167_im;
    _T_6169_re <= _T_6168_re;
    _T_6169_im <= _T_6168_im;
    _T_6170_re <= _T_6169_re;
    _T_6170_im <= _T_6169_im;
    _T_6176_re <= Switch_4_io_out1_re;
    _T_6176_im <= Switch_4_io_out1_im;
    _T_6177_re <= _T_6176_re;
    _T_6177_im <= _T_6176_im;
    _T_6178_re <= _T_6177_re;
    _T_6178_im <= _T_6177_im;
    _T_6179_re <= _T_6178_re;
    _T_6179_im <= _T_6178_im;
    _T_6180_re <= _T_6179_re;
    _T_6180_im <= _T_6179_im;
    _T_6181_re <= _T_6180_re;
    _T_6181_im <= _T_6180_im;
    _T_6182_re <= _T_6181_re;
    _T_6182_im <= _T_6181_im;
    _T_6183_re <= _T_6182_re;
    _T_6183_im <= _T_6182_im;
    _T_6184_re <= _T_6183_re;
    _T_6184_im <= _T_6183_im;
    _T_6185_re <= _T_6184_re;
    _T_6185_im <= _T_6184_im;
    _T_6186_re <= _T_6185_re;
    _T_6186_im <= _T_6185_im;
    _T_6187_re <= _T_6186_re;
    _T_6187_im <= _T_6186_im;
    _T_6188_re <= _T_6187_re;
    _T_6188_im <= _T_6187_im;
    _T_6189_re <= _T_6188_re;
    _T_6189_im <= _T_6188_im;
    _T_6190_re <= _T_6189_re;
    _T_6190_im <= _T_6189_im;
    _T_6191_re <= _T_6190_re;
    _T_6191_im <= _T_6190_im;
    _T_6192_re <= _T_6191_re;
    _T_6192_im <= _T_6191_im;
    _T_6193_re <= _T_6192_re;
    _T_6193_im <= _T_6192_im;
    _T_6194_re <= _T_6193_re;
    _T_6194_im <= _T_6193_im;
    _T_6195_re <= _T_6194_re;
    _T_6195_im <= _T_6194_im;
    _T_6196_re <= _T_6195_re;
    _T_6196_im <= _T_6195_im;
    _T_6197_re <= _T_6196_re;
    _T_6197_im <= _T_6196_im;
    _T_6198_re <= _T_6197_re;
    _T_6198_im <= _T_6197_im;
    _T_6199_re <= _T_6198_re;
    _T_6199_im <= _T_6198_im;
    _T_6200_re <= _T_6199_re;
    _T_6200_im <= _T_6199_im;
    _T_6201_re <= _T_6200_re;
    _T_6201_im <= _T_6200_im;
    _T_6202_re <= _T_6201_re;
    _T_6202_im <= _T_6201_im;
    _T_6203_re <= _T_6202_re;
    _T_6203_im <= _T_6202_im;
    _T_6204_re <= _T_6203_re;
    _T_6204_im <= _T_6203_im;
    _T_6205_re <= _T_6204_re;
    _T_6205_im <= _T_6204_im;
    _T_6206_re <= _T_6205_re;
    _T_6206_im <= _T_6205_im;
    _T_6207_re <= _T_6206_re;
    _T_6207_im <= _T_6206_im;
    _T_6208_re <= _T_6207_re;
    _T_6208_im <= _T_6207_im;
    _T_6209_re <= _T_6208_re;
    _T_6209_im <= _T_6208_im;
    _T_6210_re <= _T_6209_re;
    _T_6210_im <= _T_6209_im;
    _T_6211_re <= _T_6210_re;
    _T_6211_im <= _T_6210_im;
    _T_6212_re <= _T_6211_re;
    _T_6212_im <= _T_6211_im;
    _T_6213_re <= _T_6212_re;
    _T_6213_im <= _T_6212_im;
    _T_6214_re <= _T_6213_re;
    _T_6214_im <= _T_6213_im;
    _T_6215_re <= _T_6214_re;
    _T_6215_im <= _T_6214_im;
    _T_6216_re <= _T_6215_re;
    _T_6216_im <= _T_6215_im;
    _T_6217_re <= _T_6216_re;
    _T_6217_im <= _T_6216_im;
    _T_6218_re <= _T_6217_re;
    _T_6218_im <= _T_6217_im;
    _T_6219_re <= _T_6218_re;
    _T_6219_im <= _T_6218_im;
    _T_6220_re <= _T_6219_re;
    _T_6220_im <= _T_6219_im;
    _T_6221_re <= _T_6220_re;
    _T_6221_im <= _T_6220_im;
    _T_6222_re <= _T_6221_re;
    _T_6222_im <= _T_6221_im;
    _T_6223_re <= _T_6222_re;
    _T_6223_im <= _T_6222_im;
    _T_6224_re <= _T_6223_re;
    _T_6224_im <= _T_6223_im;
    _T_6225_re <= _T_6224_re;
    _T_6225_im <= _T_6224_im;
    _T_6226_re <= _T_6225_re;
    _T_6226_im <= _T_6225_im;
    _T_6227_re <= _T_6226_re;
    _T_6227_im <= _T_6226_im;
    _T_6228_re <= _T_6227_re;
    _T_6228_im <= _T_6227_im;
    _T_6229_re <= _T_6228_re;
    _T_6229_im <= _T_6228_im;
    _T_6230_re <= _T_6229_re;
    _T_6230_im <= _T_6229_im;
    _T_6231_re <= _T_6230_re;
    _T_6231_im <= _T_6230_im;
    _T_6232_re <= _T_6231_re;
    _T_6232_im <= _T_6231_im;
    _T_6233_re <= _T_6232_re;
    _T_6233_im <= _T_6232_im;
    _T_6234_re <= _T_6233_re;
    _T_6234_im <= _T_6233_im;
    _T_6235_re <= _T_6234_re;
    _T_6235_im <= _T_6234_im;
    _T_6236_re <= _T_6235_re;
    _T_6236_im <= _T_6235_im;
    _T_6237_re <= _T_6236_re;
    _T_6237_im <= _T_6236_im;
    _T_6238_re <= _T_6237_re;
    _T_6238_im <= _T_6237_im;
    _T_6239_re <= _T_6238_re;
    _T_6239_im <= _T_6238_im;
    _T_6242_re <= Butterfly_5_io_out2_re;
    _T_6242_im <= Butterfly_5_io_out2_im;
    _T_6243_re <= _T_6242_re;
    _T_6243_im <= _T_6242_im;
    _T_6244_re <= _T_6243_re;
    _T_6244_im <= _T_6243_im;
    _T_6245_re <= _T_6244_re;
    _T_6245_im <= _T_6244_im;
    _T_6246_re <= _T_6245_re;
    _T_6246_im <= _T_6245_im;
    _T_6247_re <= _T_6246_re;
    _T_6247_im <= _T_6246_im;
    _T_6248_re <= _T_6247_re;
    _T_6248_im <= _T_6247_im;
    _T_6249_re <= _T_6248_re;
    _T_6249_im <= _T_6248_im;
    _T_6250_re <= _T_6249_re;
    _T_6250_im <= _T_6249_im;
    _T_6251_re <= _T_6250_re;
    _T_6251_im <= _T_6250_im;
    _T_6252_re <= _T_6251_re;
    _T_6252_im <= _T_6251_im;
    _T_6253_re <= _T_6252_re;
    _T_6253_im <= _T_6252_im;
    _T_6254_re <= _T_6253_re;
    _T_6254_im <= _T_6253_im;
    _T_6255_re <= _T_6254_re;
    _T_6255_im <= _T_6254_im;
    _T_6256_re <= _T_6255_re;
    _T_6256_im <= _T_6255_im;
    _T_6257_re <= _T_6256_re;
    _T_6257_im <= _T_6256_im;
    _T_6258_re <= _T_6257_re;
    _T_6258_im <= _T_6257_im;
    _T_6259_re <= _T_6258_re;
    _T_6259_im <= _T_6258_im;
    _T_6260_re <= _T_6259_re;
    _T_6260_im <= _T_6259_im;
    _T_6261_re <= _T_6260_re;
    _T_6261_im <= _T_6260_im;
    _T_6262_re <= _T_6261_re;
    _T_6262_im <= _T_6261_im;
    _T_6263_re <= _T_6262_re;
    _T_6263_im <= _T_6262_im;
    _T_6264_re <= _T_6263_re;
    _T_6264_im <= _T_6263_im;
    _T_6265_re <= _T_6264_re;
    _T_6265_im <= _T_6264_im;
    _T_6266_re <= _T_6265_re;
    _T_6266_im <= _T_6265_im;
    _T_6267_re <= _T_6266_re;
    _T_6267_im <= _T_6266_im;
    _T_6268_re <= _T_6267_re;
    _T_6268_im <= _T_6267_im;
    _T_6269_re <= _T_6268_re;
    _T_6269_im <= _T_6268_im;
    _T_6270_re <= _T_6269_re;
    _T_6270_im <= _T_6269_im;
    _T_6271_re <= _T_6270_re;
    _T_6271_im <= _T_6270_im;
    _T_6272_re <= _T_6271_re;
    _T_6272_im <= _T_6271_im;
    _T_6273_re <= _T_6272_re;
    _T_6273_im <= _T_6272_im;
    _T_6279_re <= Switch_5_io_out1_re;
    _T_6279_im <= Switch_5_io_out1_im;
    _T_6280_re <= _T_6279_re;
    _T_6280_im <= _T_6279_im;
    _T_6281_re <= _T_6280_re;
    _T_6281_im <= _T_6280_im;
    _T_6282_re <= _T_6281_re;
    _T_6282_im <= _T_6281_im;
    _T_6283_re <= _T_6282_re;
    _T_6283_im <= _T_6282_im;
    _T_6284_re <= _T_6283_re;
    _T_6284_im <= _T_6283_im;
    _T_6285_re <= _T_6284_re;
    _T_6285_im <= _T_6284_im;
    _T_6286_re <= _T_6285_re;
    _T_6286_im <= _T_6285_im;
    _T_6287_re <= _T_6286_re;
    _T_6287_im <= _T_6286_im;
    _T_6288_re <= _T_6287_re;
    _T_6288_im <= _T_6287_im;
    _T_6289_re <= _T_6288_re;
    _T_6289_im <= _T_6288_im;
    _T_6290_re <= _T_6289_re;
    _T_6290_im <= _T_6289_im;
    _T_6291_re <= _T_6290_re;
    _T_6291_im <= _T_6290_im;
    _T_6292_re <= _T_6291_re;
    _T_6292_im <= _T_6291_im;
    _T_6293_re <= _T_6292_re;
    _T_6293_im <= _T_6292_im;
    _T_6294_re <= _T_6293_re;
    _T_6294_im <= _T_6293_im;
    _T_6295_re <= _T_6294_re;
    _T_6295_im <= _T_6294_im;
    _T_6296_re <= _T_6295_re;
    _T_6296_im <= _T_6295_im;
    _T_6297_re <= _T_6296_re;
    _T_6297_im <= _T_6296_im;
    _T_6298_re <= _T_6297_re;
    _T_6298_im <= _T_6297_im;
    _T_6299_re <= _T_6298_re;
    _T_6299_im <= _T_6298_im;
    _T_6300_re <= _T_6299_re;
    _T_6300_im <= _T_6299_im;
    _T_6301_re <= _T_6300_re;
    _T_6301_im <= _T_6300_im;
    _T_6302_re <= _T_6301_re;
    _T_6302_im <= _T_6301_im;
    _T_6303_re <= _T_6302_re;
    _T_6303_im <= _T_6302_im;
    _T_6304_re <= _T_6303_re;
    _T_6304_im <= _T_6303_im;
    _T_6305_re <= _T_6304_re;
    _T_6305_im <= _T_6304_im;
    _T_6306_re <= _T_6305_re;
    _T_6306_im <= _T_6305_im;
    _T_6307_re <= _T_6306_re;
    _T_6307_im <= _T_6306_im;
    _T_6308_re <= _T_6307_re;
    _T_6308_im <= _T_6307_im;
    _T_6309_re <= _T_6308_re;
    _T_6309_im <= _T_6308_im;
    _T_6310_re <= _T_6309_re;
    _T_6310_im <= _T_6309_im;
    _T_6313_re <= Butterfly_6_io_out2_re;
    _T_6313_im <= Butterfly_6_io_out2_im;
    _T_6314_re <= _T_6313_re;
    _T_6314_im <= _T_6313_im;
    _T_6315_re <= _T_6314_re;
    _T_6315_im <= _T_6314_im;
    _T_6316_re <= _T_6315_re;
    _T_6316_im <= _T_6315_im;
    _T_6317_re <= _T_6316_re;
    _T_6317_im <= _T_6316_im;
    _T_6318_re <= _T_6317_re;
    _T_6318_im <= _T_6317_im;
    _T_6319_re <= _T_6318_re;
    _T_6319_im <= _T_6318_im;
    _T_6320_re <= _T_6319_re;
    _T_6320_im <= _T_6319_im;
    _T_6321_re <= _T_6320_re;
    _T_6321_im <= _T_6320_im;
    _T_6322_re <= _T_6321_re;
    _T_6322_im <= _T_6321_im;
    _T_6323_re <= _T_6322_re;
    _T_6323_im <= _T_6322_im;
    _T_6324_re <= _T_6323_re;
    _T_6324_im <= _T_6323_im;
    _T_6325_re <= _T_6324_re;
    _T_6325_im <= _T_6324_im;
    _T_6326_re <= _T_6325_re;
    _T_6326_im <= _T_6325_im;
    _T_6327_re <= _T_6326_re;
    _T_6327_im <= _T_6326_im;
    _T_6328_re <= _T_6327_re;
    _T_6328_im <= _T_6327_im;
    _T_6334_re <= Switch_6_io_out1_re;
    _T_6334_im <= Switch_6_io_out1_im;
    _T_6335_re <= _T_6334_re;
    _T_6335_im <= _T_6334_im;
    _T_6336_re <= _T_6335_re;
    _T_6336_im <= _T_6335_im;
    _T_6337_re <= _T_6336_re;
    _T_6337_im <= _T_6336_im;
    _T_6338_re <= _T_6337_re;
    _T_6338_im <= _T_6337_im;
    _T_6339_re <= _T_6338_re;
    _T_6339_im <= _T_6338_im;
    _T_6340_re <= _T_6339_re;
    _T_6340_im <= _T_6339_im;
    _T_6341_re <= _T_6340_re;
    _T_6341_im <= _T_6340_im;
    _T_6342_re <= _T_6341_re;
    _T_6342_im <= _T_6341_im;
    _T_6343_re <= _T_6342_re;
    _T_6343_im <= _T_6342_im;
    _T_6344_re <= _T_6343_re;
    _T_6344_im <= _T_6343_im;
    _T_6345_re <= _T_6344_re;
    _T_6345_im <= _T_6344_im;
    _T_6346_re <= _T_6345_re;
    _T_6346_im <= _T_6345_im;
    _T_6347_re <= _T_6346_re;
    _T_6347_im <= _T_6346_im;
    _T_6348_re <= _T_6347_re;
    _T_6348_im <= _T_6347_im;
    _T_6349_re <= _T_6348_re;
    _T_6349_im <= _T_6348_im;
    _T_6352_re <= Butterfly_7_io_out2_re;
    _T_6352_im <= Butterfly_7_io_out2_im;
    _T_6353_re <= _T_6352_re;
    _T_6353_im <= _T_6352_im;
    _T_6354_re <= _T_6353_re;
    _T_6354_im <= _T_6353_im;
    _T_6355_re <= _T_6354_re;
    _T_6355_im <= _T_6354_im;
    _T_6356_re <= _T_6355_re;
    _T_6356_im <= _T_6355_im;
    _T_6357_re <= _T_6356_re;
    _T_6357_im <= _T_6356_im;
    _T_6358_re <= _T_6357_re;
    _T_6358_im <= _T_6357_im;
    _T_6359_re <= _T_6358_re;
    _T_6359_im <= _T_6358_im;
    _T_6365_re <= Switch_7_io_out1_re;
    _T_6365_im <= Switch_7_io_out1_im;
    _T_6366_re <= _T_6365_re;
    _T_6366_im <= _T_6365_im;
    _T_6367_re <= _T_6366_re;
    _T_6367_im <= _T_6366_im;
    _T_6368_re <= _T_6367_re;
    _T_6368_im <= _T_6367_im;
    _T_6369_re <= _T_6368_re;
    _T_6369_im <= _T_6368_im;
    _T_6370_re <= _T_6369_re;
    _T_6370_im <= _T_6369_im;
    _T_6371_re <= _T_6370_re;
    _T_6371_im <= _T_6370_im;
    _T_6372_re <= _T_6371_re;
    _T_6372_im <= _T_6371_im;
    _T_6375_re <= Butterfly_8_io_out2_re;
    _T_6375_im <= Butterfly_8_io_out2_im;
    _T_6376_re <= _T_6375_re;
    _T_6376_im <= _T_6375_im;
    _T_6377_re <= _T_6376_re;
    _T_6377_im <= _T_6376_im;
    _T_6378_re <= _T_6377_re;
    _T_6378_im <= _T_6377_im;
    _T_6384_re <= Switch_8_io_out1_re;
    _T_6384_im <= Switch_8_io_out1_im;
    _T_6385_re <= _T_6384_re;
    _T_6385_im <= _T_6384_im;
    _T_6386_re <= _T_6385_re;
    _T_6386_im <= _T_6385_im;
    _T_6387_re <= _T_6386_re;
    _T_6387_im <= _T_6386_im;
    _T_6390_re <= Butterfly_9_io_out2_re;
    _T_6390_im <= Butterfly_9_io_out2_im;
    _T_6391_re <= _T_6390_re;
    _T_6391_im <= _T_6390_im;
    _T_6397_re <= Switch_9_io_out1_re;
    _T_6397_im <= Switch_9_io_out1_im;
    _T_6398_re <= _T_6397_re;
    _T_6398_im <= _T_6397_im;
    _T_6401_re <= Butterfly_10_io_out2_re;
    _T_6401_im <= Butterfly_10_io_out2_im;
    out1D1_re <= Switch_10_io_out1_re;
    out1D1_im <= Switch_10_io_out1_im;
    _T_6402_re <= ComplexAdd_io_res_re;
    _T_6402_im <= ComplexAdd_io_res_im;
    _T_6403_re <= ComplexSub_io_res_re;
    _T_6403_im <= ComplexSub_io_res_im;
  end
endmodule
